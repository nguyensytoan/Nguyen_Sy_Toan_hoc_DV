// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
e+Kh9RAQTc1VGgtdAwh+d425Ebn3MPduUsJaKtfDLxs3qcwMefSl2azGSOo/sMbNtnwalOVVUNsG
eDgndbfMWIyB44MnBRfIxkcG9wStN/Hb9qwzghs/xN//XokpmCkO6JacqTR+x0pQbzR9Obrpeq2h
dIJ3hlpJiZ4l3rqZTLHDX8k1aiMNaS9heNEMwTHKiO6tGLOmNcuY5DQket5kJvw8/+96/qNherCk
+DVYVfQD7Db34ByxBLQzmHbkUmCMTXfIm4Fc+dcSG3pNY+BIIzRqm9v4VYDcZ2L8RooAQxFuLhvW
N7i/Rqvu/KqAFJwz+lwXQ6nC22Y3f0OxC2Nmew==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 12352)
NoOWvFZrlR7G6IjlWB5J4j7ZuKeC6gzRs2sLKmso/QKyHUUYMW8ff0VrljLKhki0t3Tpq6Vg5lYS
l9GSV5Fy/Y3/67aPEmK3c9SbHGS8uT6mb/oF2dPYx8igqGNBJrVSWIQ0nni7xGkOamq+5FCWsalY
9wxs4g+j7pJQNkBRpHJPj7JP4Rzv4sr9d4wCeVi0EZb5O5VAZS6pvFzgGo+kgAsuJ0iIjr59/7IH
fco4UN4GhhLBZdz2inoMDfGpRjp0i3NQqsepmLoaSxp8tLH3TpFpQqx1xMnN3PHORavP7Jwi9yDs
js7ONoZDzUx7KtBZeCPe8v/xzW25ENdULy5QN8A6jtwPXf+FAhF44vbW85Ql12Z1EIm32wIML5FJ
8sqVadl+xg7vozw+dEszGCR42F5CAQi0TF1dW7xk/b77S2qBnYwsW5q2I9HmSgII+7z+LVMcE15b
5Dmf8t+bxrMf7kuvyl1+OrAbNkrjBZ555OacwRz/mLrwTfc0ynUv7pvDD1tihy9QaBH0z/+rs/OQ
Hm4qlYptL43alAWXW09ZVrtqxPDhz9zk4iKBiDG/R+fkh7G6eCnktwD3/H19LabAg1Zx719F1Xn8
4KiVQgOYdJAMJGASEnaVs/fhywZlV3FYH84t66V/QbRmlkuxGL86tkgeHSFtiMnd1Mop0ZDWoRgz
dx1GSiQHwppLqI+ZSmrhC7Tjv5NkIgy6nNCE0AVkM2skpDVQZh/UtWpy/3d+nblSK2VCvdrhyI+D
qps3H4CpVSIHeHk5SSSzsRdQGWDA0FdkclPMok9wLtIpY4CZZmUsxu/nGBfKIOB1OUFsnxRm07j0
zc5PFDfgYyX8KdPLX/iPD1bsFL3ew3V5q86J8WBEmZLDmJhfrcfa42G/r6J55up4wKTtoqS6qQUu
l3SNoV0+1fizmU+v3+ilrvb5X4aP5uUdnEvqjooQPgQDz+fOt2y879q6HWF+VyY8D0RuPef5PPco
mLUt1i09UDK14ldz8jTqFBAIum4RmB2SSOrhG331GFZEZQXTwqvF1Q+VnDxfy5tpyCe+3ldo4GHu
s/lHoMYpfBKr5mMeKP/rylKU0al2+emxVp7MTUo6ie3u9CB1KnndmdmxDcUuJgD+BDCaMRBBHu3c
Cma1y6hy3Yt9QP8BZcT7ZY1L9Ej32hJL8a2rqYdHUJ25TqpkTyhmoJjX1UySMhKCgi2QrDH81JFH
PGzD3YYk3PqVNxzkCM7pWaY2icVzD3RppWNSmXsNpmRxUL6IPldTr/xXHy3vK99ASeom+mPJBKfw
/+oWmaZOl6FmKJImXwCYBgJUlPHlSkisFKQlKmOnluMwUsYnT/htcgcTiUY5Ipc1liE6QXMU3Ox0
8KpI+f6QjVtdqsQqU17+2asNFuKHe39tpyfXJZpOFmaIa5408Q/BpCCuhvu/pHEeCiaepYo05iQm
5ssiEEF0s03TTK+s+6WaE3BWPgizGuQSc7Tvh9hBDH8LkSQYynWsJ1Dq/RtztCik1q72W9bKblOd
/wOQ0JBqgdC02eJUQCc6HfQiXo4oTKnfl50FQ5S4doi1OTFazJva7FFEhnh8fb6B92PKPJAzYoUJ
2Y77Pqo3cr4pao0SqaSN8ZpURhYO/VujZQS3zfQ3c7XDftSrpmIMdyoDB0vXgnZ4xEE+dntWxdSZ
6k4JPJV2bgVduoiEH4YL9ImBiGsdQcNrqH2dl+wo3sr1yRG4mZY/ptw3+Pmd6/ZvjqyxcN+Q5MDE
nehFTz/wrtIAWZTg+s8slkLJ33VqWX9up/PTU0QgoUJrRVU+1e8TosSbZ2xjEXhb6XDSUgZO8Ick
RIDPTpb5WtskFvs0mBKunYiLr1mUdLE8gsoycrhnnKxijvozJabIiQBwFL0QRMlvgbMhV2dWIXtw
yqjHd+sEi5Up8xayoQBGjkdGip2qUE7p5gD/eiEdbs0ozo97bKW9S41jidJ957c0njWwhGjh6c63
+Lqfh9Dh5UprlCF5vptqlvGOelDE6f36dRscB0bsDVHNAmbtbWu1kyz0OYpz2xSgTcUhFDIOQbKr
bXPFTANNQ+Sd9FPRRuCYJkI8aZ59BlNj2kxUAjBKfmhA74fucDnP1nbzz6PFw4wcLCU+eLC6BzpH
WLAPGRMlcjnw7JlBoqkizK1l8cBcFCkW1kOlLv4bnuD0PHpIPOrKgq3GTGJnkqwq5mTDQ+Oe4dGL
cl3k+uI+52o7H71c34BqGcCD9s5InHbEyOGzBR/Y9W82NedMQ+YlrawTixkoIKyaKiW5+ew/gtT2
Z8FHrLKfDlVKEYuFAUGJgN6d5vT8i9aNqzFMHBWnmz+7K5tCaGKsNINl0RCZW5QrIrM/CQhggwD4
r1dUKw5ZGH2SDWKCRcsEIjhrR0ffDvKVWWSsRDna+keviwjeag190j2le1PekEIg5iHrBhpxNECk
dyt+VfNVuE5laIqAEFHMiGb+kJ+jV0FpSf+a7CE+uQo1HeY4ap5EzgXGu68Mgp4BTmX0afAwSsbq
9g4x36IhZFk0TmKETh3Opno3n4dknNtUe/KBWBWtZwQnOZ2B991hcAQVXLQ5DNHDE8vNy43RJwux
s4eYcr6rfyMDE7DJGmBx/JqO1dH9lacUxmjRmtzM+5JoFAMexMwHfJf/G0+GLSTMKEd4BviX+OKX
Bu7p0MHl6sIQ4Uu7RUhTAy4eEm1tWvONiAvVkFHbII/++cbqr2j0+7iBBQXP6dmL6fEpFgNaWpP4
dQ17ewNZm2YQZggjBulcASHTnS7rDM5VMe/1Ta42ZRhN6TxbLtq78vsW2J3zoSIQTgSvg0NBgokc
K/l4HkQnalQp1E6nsl+4nFw8tXfJmOH34QC4GAolTy4jOugFzF58K8nl/hjM7phQrXjqN4l+s6g2
ZYgch0n1Opsk6cNMhIaa261X2/r4ajIzcLsSmmUuxfERKpmirlk6Qy5HbUQSU3B79OoAua4Ca2zd
HWvtAHu+kx5W4Pyw6teeH9x7G/IgUC/iPt/S6Y4u3WKqlf0EWBaa8xV8iVEW3M2fwtYpd8Z05pD+
GXNz8TIBTT418pdy6+2IWCwa8ZS4cxPHuwLOEUM4IKSc+gnSCT1hoM+VlxW7xZdKA9TNz24y1m/Y
596osIwueVkfowzUEZV/GwZfWDRS5qZjMyN05FLFkEZSEeyBp7B263H6D2hkhcJaNHt8KL/wixDt
Tv8D+oeuwvbHm04xmv/DxPRPwIT1sSXWQPwevPje9pOQpOq0ciDHNq/zBf6EmA1wQzcf9FEG68kt
MJ43r9IWxtG+dVGCX5oClQh+TQIPs/ihpq5VJx29KNThmFgGJKrng06UWiHtVE5IKlYdnD4welmH
C71C7y1GrjVtWZsXVWIbRX4ipc5l3kG/l6AYxxjw3SVhn9ryFEUZFa16eyj/NT8uM/C04IVBpesM
9zo9ZgqptisvKgzm0BjRhY7xfUDRlWTlC71PTa+H7IbfPtmq0bS7eVrY6sHXktFeAs5ZRh13mtaJ
JnDWI6tJ9MlxKTjabqzXfh1EFP63CvwQLTyrn+SQ0n0wcdjYBzaO4XuLF7jbhzm+ZtACw9Hfq+f9
zSqe9Aic7PyFopwC2LU5Y4d1uiHyzdxuJolk1F23+M+QWrdPRtq5icHKEhA/F0sp2PBSusfijpFO
+MAUuES4ZnzQseGd2iBF93BQmjlm2RxzEV5fpdOR2aVmZjkakxQJWu6URt5wmPom1gjs8pcvYz1A
EHXntCCUpqE/YBAjHigQeT2/UDINMwWgKaL3GFd9y/FYjUVHiw9SEr88V2BdhaU/GyCrQUuQE5zw
1CI6APYFPYxp+XYoFjMZ8bhEWpp+KGNnQ8EosMer3GSktMY8Xc64eY1aPS2ijXP/VRcNGzWpsNrc
NFuzbtxdKoYHNGZm4lLhWcrt738/vgbsnVsJq3LORKexNNsXWOIKL1fhCClFMhYPNIswenLz1CXc
pnBD8u/CWC/f8h8/XUHT+i3njQT2OXzoPPq2e9sY2lIh+1dDsf1sJ+8wz6j+I+mQQWuzdu1P6CH5
MfRBSsGHPQU2kr4vJD7gWfi7dXoFM5eGBlTwSLq4ncFrm59v5Lvp+0Vyt8Op54DYQjeJ/pAT/WpK
S4RRJ0GD1nm0FuJjWTHEKCiUB5sDqz8Ft5B7tCRV7vLlY+waex3OYLXqLtBSnp1hb5qeD/fWGBpK
2ETO6Ya9lziQ4WDkF2KKms7rp9D4Ctzw2unfOKrOv3ldyK1ivZbWTKMAtof+7xR/V/nK4/OMenYe
QhT0oC080Kn0cu7S0ZDV7P4t2FeXTYcATUAFk7Lh5xB/fefWLT1+RpfJ3GH4rBj6Qqkr35Fu6HAN
CDGMumnuF/yZv6YgIC2nGHSqSN/nP4/VQeJqOmnStTtmoNkxn5IkbNs85akVTOCbxwr+a7NIcjUP
IyAiVDOJ+5dhlvMI1q9ivq10c6mb2w8ZF/mwvFRWBCNYUi/ixpgb/vDKuhMGld7bSLcNtVglPkUe
IeCH7ASHlnOT23m7rJNl5Wo7PcePa1At7Nl7NMFvG57XISf0vzhlAnfP/roQBJ09pm2INfJ3R4cv
UchrEqZkuhDNGxbK0VEFMvr3E0GL/jVCcvfjLpUS+IVyA4gAYTXRoCs0E72edmKipnwQ76vhSJIK
nVVkpe3uDv89en5bGwNutldMob7iFX9O9VgCosovqaDw0HaLcMpF25p+J2f8lT/xRPRaYUIeW66C
sKSvwKLN+EKHTYX65VcMi1B2OAr6b5P5W/RikpYa0i4lGQwM7IF1NJSF7r/zKP9lfTnE0htSDeJ/
z7xe+ENH9YX+emKy8kH8bKoYDp074RdgmtYajh2Axrq4qZ+TD4W59ZeCPnUlN/y7HbSQrPrmmvYH
uJFRu0PRUU2ABOQo7nB+KCQAcfTs6xmsNa5QOrDRM+B1Wz9BnEdwvH7h3LsVa+x4NCN2CHbdiuc+
hhbzQ5yFKQGZsGD09zqB0wJo+Vpz7n1hNIqD39cA49eaOMhC878KGKf8I2+YQXok73VK6juOz/kO
orvsOEy+XIYl9aOSUk4gqxO5wDtkvCEalaveYsyG5WIRJ403Nftb5z8uEMjW8fWPmeoQ+26TkUMV
5UHX4kZNQ39+FBFF4mpFuURm+d6c6p/0F7/rpBuMSfXH65AFh0SvBfBQPRQJ9NQwAuGiBbuKl8Pr
luCOaKykbBFP76P8yv8WjZFxuuqNip8B1hB3IT0gWAKa1o0R1n0a1TAp/+LHcTZbSfdRlWBPasB6
8sk3VwRfmoujqaR3MrrPU6eUlDgBIbuy30weAx3e9KIXKaHb/dp1PaIPLQeSvuSjkr8FTi9NCdCR
WvWmFaHvdQ3a1hQpaiqNpHVVerdkI+31/byEhEGd6HgdvuQjhrwRgXtMpimxX/pTRVtKZ2nLp7+G
tcB2Me5mfEM1MHAHaIxEx9yrp8LUp08QCqa8h19xPfGd0RLL8qHPMw9atB+eX33P4pIcG62NBlce
vUJh2Sj5PPoReqfLCe4Rx41EhfFkqvPvr99bvI8bRvCyU8Hw3Z4thCbLdC+wUZp2nRI9DYOuVKot
NjluLfxFPrIr92Bkc2v55fmp6KG9yX5nH++SAJWggYVJaDUrzXBakNt0xM5x/4tT+PnpKzy9qgkl
U7N6Jb3VWt7GSy4PZSlnyEok3TBFZty75ryQmTG6l1qdmOrCoCfIUWNDI3QSi08B3wKuvIXPaKiv
QZ0lidXBiji7HKe7g4gx9shYLd9Px6AJG148Kd+iUoSohbrZr8TAqdkdVyomZtIB2iIVIUMbLA66
ADOHieZG1upIfvgJ5AvNtyitFRB9KjR1PoHKw0Y6WdaZxIyziRnIDGC4DilLfiwY2GTgCuNw0LS6
+t8XxTJKkbSRsakE0dkne0jhbjnZ6qilZ8dLnU7ixlgy5gRGecPJFjA8myjMeH2Me0ICj1BfzyrJ
jXd5qdyVG0GbqckiB+BM8qVLCs7M/ZI43HS2wYLBMXlXsemH2Y6fdmCnUIPupkTeGyylcpG9c3sT
WMs9L7G9qpwbqPUo2Sl5Tnwbn5SZ96CWCmusnKHqIYzAXGdvUdz+0E8XyEK7qFVT5NqqvDw7zehO
QnaYfxYZyUei/mDLkC1isx6xSSe6PeR/Qcz4Nn6ethF0YlCxHLea3Dk1mllmcigVPpNB85rXRoSz
dWdMOFkBlxICYyHMK38QVuknWmyzj1Kt0RsruQFcao28vk8HXb9hcU+yBixFpnXtvsel9xSr4Ifa
H0iiBbo80UnCb/SDeWyZZpU8ifzT/SzcI95uXeyoG9cVSVNBp/F8lpidC1AbkERTiyIpdY3BWZoi
FVfUwiN/dRYn9XX7acguBZLn2E7tbtAOSkWQblNM85cp6k3wNxC5iCkRWXpKEzNcp46v4myrRhwL
q96Yqrg+0xmnHRusrBZTuAAjLLAWACrrqrJCbKsuT3b+KCTAIzujlNbw/U5m5K/cbF0aL7rUMYYq
4pjUzpCFG1eMvL799AqXpNIrScQVuiHVuBD4HK+TKQ2couGEc1Qz83anKqGIf24BBCfxxPlRccqL
y39BI/FFSVkZkwHeji2IwgbgsyCGwHEAjruriRrXT8loktB3LzYoV7TnFs6/AT7D7wRuy3VW++uT
uJciUIitnjHVC8wFFuunCpTL2Q5jTr9UCRfmPfvqaEfn+KFyzH0SJtKK5eT9H7BIm3Mq6uHFsdfs
OiwIljAKyVu1wXOP0FbLy9XTm9iBX/DhIjrBlCzpb7bip9yTukr00Ji68fwKv0GD9EVntGKm9Zmt
UPFS+Von1uFi0UrNLXC1lO4OrL0wAFxrY9ynLxI4EWQZ2oFkksdDXW29BWrKVLmzs2ns3pRrzVaH
keZz/fkkJEo+gLTlw77Kyy4kGZD2qqecBI8JpcjkQbe3ts8ApaSE1GkqDUHmXqOzoOtYgedOErkY
zhwdtztQSSOOcys9LPRlrpy5TupdmnZb8U9ktCu6Su9wFdFAIlouyMetjy55/SiVz9ZYfZpR8SIf
M2BDJ9pZW4xZJyQstUN9tOTSgMIv/V8EwcLdvpuDwGcPAruM3/66FwlQS5aeqW2uI9/n+tmMCPqU
6dPIpvDdUCwI7MuP48JzxzMSKs/sxYdsnapo25cUPi4IyzZDDjG6xZ4pWHyCCPJnjCJzOAWuyher
sz+Zu+EIgtVfcOMLAQpGy+Q4yXcd6PVyo8fgC/gi2dI5Nx8zTt53lnffkxxwO0Jl4s1ALdZBDWOV
/DDdDLgDpatxzMFOtB7pt48XFjcBJ96ypA8GpMSOf0yNqqFRsN5G8iu5C60qrlicEctydt5kML6I
Ml1R0ae1aWHHRLFJv6W3GiosnYumkdY3N7RA8gSkbgF+vDjwvY6tUOUM6aOvrWFOuuPIeaPR/Xec
vjVboZkmxTdfWqZbJJDR4Ht2lXsPtuHs/vUoqVJhbA3vf8eXRwENGvrV8tS9ZPVNbLGPib0CqyZB
Y1ReVJEjYyi/2rAM1x16zcFPpR4nn7mdXD91+kYynz4jmJjq5K34bphO1KDSfvAeQu5fxBPfXsYg
cosAg/zqXGTikwFE1wWyfjG1Yc9cj8XEyq7or6PrkxSR1/pDUNvAEPgjN6LByPyw85Vlr64eqpvO
+DoBkZFBrQ6HxmpEnAahvHXyQbXmrhomcVda5h38p+7wgTXvgQPXImVVImMuIHcKE5GNQg/FvPY7
5sQpZZZ4bSzOuulMUI9JGLdI77BxMCNYgm1Up/XCWSAU97S8foVE3jLIHy2+lWwCbNXBz9owg2eP
G0z0gZqA+/+ZwKFKJ6ZXdQnnNHCbcnBYwHGqZ9sPPtAZtfvNGOVg8RgjXre9P1xz1Omj5gsU4URH
LaCfFWBsNPmTc0p5thD28QcPcbydARBfZ+NWytzuTIpYXVu6pahJSKEx0n6vUGkrd7ms6XIxfLHA
Xod/xnzA5qm2Jxp10Fq8XpsI2RIsZxLmSV2t3gER3os4iF9oZ5jAQWNY9wb9sHROPg2pKZkQyGX4
b+TKHE9UaZKdQUoPUVbcF+N3fFoe+AaFxmXrMzXINOtfMjlXGhZS92smS6XDtxesSEKC6UPy+vME
XFzvu1qk66v1Z9eaDEoHDu/gE+Th0sybvr5DspfbCcF6MfgJjOTuvchr7btADk+xOB2fZGx+He/Y
uymUILzCW1po9G8gGppAh9y6yIwwqLWpjm2NAeVfEWU3ayPfc7v2q/fRPJDntJb4JCJpDLxmR5B2
n9GMAoI7jjsWMGZ65GrFpDZNLJI8M0EhP0kMhniaL7FMTIsVxjUc1D9cZL4VX1VIk8RoVAtWkCvS
Oa3zOCWudVXfgA+GwGZkRQycAq1mdaGc8FGR+JiAYqItHcx1sKY3Ld7XNuyE4cROFRTLhGJYeFOS
5AKQv+MQGjYTC/kCPeXJ+2YSluDpSl4UFJAQdHbfrd7keIjFTvxfzfklDsJ0FrZAeNJ8AZaAtTwR
/iscAIhhjIvq5PWsWGMbKfH9cWVRNX5euBmHRp73jIdwIbML/crOyz3JkNagGiN30YNH4vwkR45H
F8woIMWTtrwT/5oDTcyFpx+P5tk2ix59DIfDUXX+GPfhJIsWpQsotddBuKDgnMiPCEV4mf3N/R5V
RUYP9Ah7zUJ3Z0zSmu2xcBzbWs1u5ShtNcdtFL0HWrh9qJMxOQP8DQbrzYFdN9DmJa5Nb+S/pSH4
xwUZl2nkBQi9hIBzVkxg/6Ll0bzQvF7Fs/RH7efP/TnRLKtsIToCRck9jJRV+LCiMghgFXjNZNfP
+Dh7cYusMIVqiiCIuU3dRhZ2vJY2IaRg65XLlx4i+fwzjPZjFDE9NVMvBYKbh5CLYzMcq/JMHYJI
GZMFk37RYd5o/kik5w4qsK2taguc8PAcE3pk6yPSSzOpDJzTa/dYo0tmv7XPq/ZzrldCDvbPrIJw
+HAix1q+9UYIxWbww1HoGgNjiK32m4CUcxoqhDWiIwWbNCQSUwpgXOpnOPt+pFrIAHTv4U5rByGJ
s4XoDUUH7DuBZbE+d1ujWrZA57BWCUQ3BPLTan1Ey8uRGbfzBHCklDyDvatB53E/+eKFWrG01vRy
i2xiwH5WUUBYpq0bhbcdWgiTeLu7BfAVBlyHuQvaUPDgwU2tYZiBi30ISjBanNl3B428U1E57lLj
gur4hl3arrOpz9djHrcaLtCpylCh3SwGGuYIfV4TWa5+5+Tkf23krOZgctQTIrL7pNCTk1FrIGKb
5kGOURR5qwovVOuOT46F1x7tat1kYjr91whLHu5LB1GieavdaPYj+yWJqCMUqSz8Zla3gVafjLa3
MITmJcvXsJVJSFFAcDBR7XUpNygscqbN5cRxwBSLZqb/qa1al3dLvYH2U1AMhzLMeZsmZHNdBv5P
kJWPtvDK6LGzH00Xamwbs2Oc8borY8EjB4QileyOYdjtcA8kFRF2RV0vbwq/6SYz5jJihG2irXxB
rIsw/5D+ivMxM1vkwyYlreTKqnYTKlmm1vkGyiPshCoRQ+dofD7ksrz8MVX3OIyvn3kTUXAj/gYd
uSgVCRe5FxBdx7CfsQkPDHSCTPHsuh8xoURGDjnomrhWpQhezD4ChfauNM1nHT48/JDeraRV6UpW
wAnTphFl4uFFuy/WsemsLwfyiuKtP1sPOdNvbpKf6xsc91nnUhMM2nXogO4802duMmLsSlyVZk3x
eqTNZPUWfpS/fqYVybNR39CQpkGzv0iyejhi4LOzMXfvd6bFaNi3r7d+a77YG0t6j5ONniAl7ftI
J5PU825LnoqaxA2LpzY5y7QlJ2xqXjCI24yTp6E7OYJvZ2R9FPtjYEQY2pFpc0BSSN3YkrEmTHyJ
RQ0SzSl4sxZ7ZBTxSxebU24xEZLXRupqNG6eWrfPL9v+cOYlQBti398gIpWm6YkH6nTG2BnVp6NP
43EPbI7oyyg9I46+Tk3kFmRaL0t1DB0n2NKG1VlmdK+0rLQDvCj8ViDc6+vzsVs83BebV7RQCe2+
OmR9zwnz2KDqkXn2+ouhx1de0RFVij2N2x/zPasr6rfygjizcg1Z8n9D/bu/wfNBMUNHErzyy0M9
7uic2DtI0fS994zCqG40AuBgCWsmalQOBcYprchQHL6antUBa/JBqyvf2phg/eXGm8iODE/+H3MT
vnEfZtqcYpHmWDfLdG64qp5C0dLVQ5VEu6CFxlInVfc36oZ5u9jFUBe2iDTzK9jxmdi2IQsdQ28b
Vgy2x7noiWOAup3GFYt/V3esPD7g4IH0SuuFt+RxGZRWMMLNHyiRqjbgEFWblsygifi7rH9NhAB4
v2GrjK5aYZEhYRSrC1or7MDDWdHfjI+qp54cAhUrdFLyNITkp5AqgtiY/NJiiKMCtPdnQNAAX2bV
pAbVI9rR8OSXDX+yX1ianqdZf4GaZDrd3LRoYxPbh1V3ICkuMy9TZAYZ22rMErKcvlIkYjSi0exI
Y8dWK7FglnOxpB4XhVQomJLqJnwh263UqZmBLlbitrp6S0oSPRoz53Z4U1HuljK20F7Tu6DpFK4e
gZtUvsZG7dyuHf9/k+gIpRI9RIaCuM0prNUh5I079feJLtf23ZT5Fq8/RNdcJXq64q+40ynGrtVq
v3oMbqoEfown0L79PpmmFUqZM2Y05c4Ud5h8q2lY5E9JWcLqgzzmoZ5SnhjDiETN7I0PN/dmi002
VHStN49k4tKBEx4ovLLqTrIStxx/AQhQ+yEjtF4MKuZtqdpqwqphSbquKFy85aRqXTs7UizFUKfZ
pNjomstQLkWBkMC7IyztCIaKRLLcUNUZQ5qlIuJV3XjSyAV6uo/EhBG8arxFugHHdS+tKJaeB53g
VW17Zp6YZM3vDzITggsSBdWjLtRf5TbO+uuEvZdFgfIK1ztfFuJTNGVb9zOP7LUVEsBRwcEvQ41E
Gf8KJKQn8fkGTEuaoXo13y5gC2BbmfRfVRpHcv+kqtvRCCawHABCoOdeHnat2n/5ie7QmEKiU8es
gc9icxyeLsJh46+p+5WBiY/ZX8L+mPSZyomB33g1iSjw0cEEdCJzNMGtdZ79Se2IYl1sPn3Qnc5u
Ksc3/Y6nJwXjN1t58Dfm38YprgP6o8/9M2tXze4GgQDG+dmQJ2wIwFRBjmXkBEtbFx6tPZdAEbvr
4cR1ntDSaTk5CJc3rp2TgzHl43NjkHnOslPPFh6c/FMZdEtdZUA1RujLnEthVOw/2rl7NTX8YAEA
14bghdoXeWS5CMKUUWpMyURhtjxSObZqg4BtvQnbfyWGEAInN0iMOJxAVKo+wgWuffnz9Ht6lWtk
K1A/kVAwbdbrphT+InU1+S4l4dwne52gq/f7tcX+pTz5C5TwYjEUjNT2cnBHezLJExEz1LY856rW
P1c0baTlS75zPVSIVw550sXo5pZCz7W18v1yvmQJuQTnWBw5MByUqYGX4S2yHaFW25WxcDv2uooi
j5MKAzeVJfJ+Kz2UR8kDyjZxO8s7i5VGFTBffXFzKMtobOqndgr6PxeVAHnAC3XA/f2rjZCwYFST
nUeTDukbt7uL2WkpDumGhe5/Wwtfos1TSbw2Wmtz9yZUOR5SH8BCIimGRZiu2AsMZs4AnDiBjgml
TeXte338sLjYVY5SnoKtwlitujmHjH2haOk5K7y0vakEVVWmkEMLKAMKCPJM11J6LXDLUFfW8NQ3
jGPS6kSKkqMH2kzowKCI5h5JrjnoEjhdkVdSwnDxbxvRR5yykhdtTmZOF/QstG8vAulcGS2CoXdN
O5ru1LCfdl5dkD1JxKgl86CdvvV9YsUEalqu0RgNCMM10/s6feIqb07fiHNiW0IVjHKOghqK2CTd
SglTIC70MEZM0XBAUwpesQc/cJjTMqGTztIiaTRpU2BAtxCRaoi4hOC3TnkMl4sJtFXwrUp5fmfC
NxP69l9j7zRbUwLKVbQSti5JjMHqi27CNHDz9l5BoAnbKbugqAoL3hrYddbtAAdOvCsIooYyW4Tp
WzQSkaRwMVwHSIbt9HHtkBqqSSyOXY+p715iEE/e+Ean921avQ551BFpSoRjaHPhFvAksRT2kiHf
kWge6yPrFG9zJAYNX5juEEIpYsDn1pm2zxmYNWfCjcPKqYCaYIPiL3D2+ptKpnjA5Nri6mhsIGSu
xlxu71+sWfgg94GJmpUC0TAsXET3qz7TOy63Ii1a9Rei4clkYVY9rqbWTdqUMJ63wfSjorJmdsaV
PKBVFRl4lP/R1msoIL51jOte5OlVRnFqtcthj1QwmmlO3SVgPfxLrPQs47IjQth5FlRUqYcCqtjG
SO02sJnTyCPQ38WvLAIzXx+cHyqT+TtuI9QZ3cwR/4PdQnSqdjAg/w9fe/a+7nw8K5FNtFfAtEWt
xCvxke0NuvRUyVlLpPZBNcG+Ay5iyqKUesvrNSHjR9vM+0CkxmwtAxU1r/FFrGlmJbHO5u3gY2U5
Q94iGNJsfd/fGQn7h/XbKvTl9D0HOC9Kns/jIJRJhuz1VNRkrb7LSM4fePEjGbxYNGoNm1CIPfvI
lse1ovp2XWMGsVLkgqcBWgD0F3XDQEkDbngVvPxae+TuWcbJnN0pVhnDuS9E6KQ8YCKGMW3omIdU
GAR3fTlSr5iFxW+dOscj0py0jy5htQxFYCmiVDbMp81zeLOQAfYxDoP1S5CVwAAKzREkeo7q+dMs
DIy5rMBIi/rgUjBWaE3hRHkcjU5+5FUoN8W5jQ5voXKw7jL4SmqXf0yq5jw6zGSwlip5uIs7dZ8c
gtCfBQk/5knNTJFb1dp71gI0dyBEUuvvVcsupXftTqe30MtsPo+KNGJxFK+9BQtBv34wRKcBWDWD
ZGSPp5TEPs3BQ3v++MaVnG+0bHWwdW+fRnjITdHWHPJ8jfAzri2z7APNCpO+3fc0D7Q7znkk6cNR
NkSxghAHC/6pgGcqwUYhW+x+aDHKVfxMj5aq+LWFbQ4kcCMJJh7TqXwbji+ZXs/F8hy+/bzqh8Nk
VdA2q4tZHoyZm4MhSsGRVzV55HZ+s/WcaNH6IycM52mUNO+1W0ILu85ei+ZdGCI0mALSueU+PUqD
XL2tjNtbF67ymgE4bv9tkELdZt7AQGaudVxS9l5ZIn4BfD9McPa9ssH5833/0kTEo/+pVNoWlzHL
IlvG7IEYytsz9I/AFWJ+UY8L7AwEnZflWpllwSKv09Hkug8Ej8FcmmIb5WBZhwCBTUi+BizgHg/f
g/mmlMpiU/ni+G5H5td1go5rfVWfp2Zx6dHRJJIXPoh4yvfdTPa1YfJXuL3KFLlQdBWkzoVAE3QP
zVYY3OYqOI8Ji+pkjkTzMSbJ0ONfeuUeEbzBgBXOB3hMw0p2g39TH5pOQfr7RFxZS5y6FmHFgk9P
3OMByH07djWhgghTdSrwSm50uwUMUVxWZVoWA1tSlSmKfblUlI60wANhhQ5Yts9AZKhoFVXpO4D3
9gf+F/X8ANNIWViYmA9d69ysjNywLWiHVBf9maCLpnv91Onec7aensRkQo0gB1hyOwLKCYX/+C1P
3BW2qsaHytv+QAgnxszDdFQyTxUMc1FxmHU+qyN4umVeapzNIkZGxYLqTmHijT2pqSGwdRVWu1gM
rLKfcDwW72D+foOCKIVGkkVNOxvtIeX0QZ3o2t7fUAFljhVn5pAaz8EaiFfEMOSaAFD9Gn0oybe7
/0l6fx5/7pf9NN/GDTNnDWdpZ8MgNxpWPmKrbD2PZxdRyIhUe4QHdZjOd+oUGgFj478OXQna2maT
PkvY0PTFPCKFWju6Np2xFyw1jlvqqS10VQMhw8IL+klx0/1aZ+PA837mZ/Kzmgx8QvJD4Zgk++Kj
TPYFLyDT7KaQlaQs36uQXOML/3Oj4GsdVP9oUPDJ8FqUnDjsr3Bvkg1LiQDHRPPIj1PfKsz1qnEU
gVrohEdH5ugRQYN3ZkPp1fvitb158dwlac4SIooNe8qv309HhrrwxAyJEfUkKu5f5RWb/jb95hy0
NYrFGheJk7ZOdZ+lZOcEPrcpEw7XUI+YVqJ3GCgLQqzysXvRWWvjFCejEMpdUjWQEjagiWatlF+W
Y2E9elV9TSqAYaZVMPxUI3sxIzfvhAuMvWKqi9rWGDNfLQxWWX6jpMjczYxi/DILQb5P+HLm7hH2
qGzBgjE93eUn8Hv0ncjHScZ/8l9oKW5fIDdUoHuxtS7NV+99HOSaO4FX84Mqh1CNa0Zw+pKbkJ1p
8EXztP5C4/51Ig6U7KGVQKqUoU8B0ZfK94zyNok5poBs6gzPSNiUfR6qr+Ld3bNoWh/SpB1q8K7+
FQbjAJpsYxZPSx+1XHvSiEKKfxvQIfeyrLtnSTaUE06M0LXOElpkZQ4P731Ip92Zup4U+3g0ypv3
Tyj98SUFuhAw2i3YnQp1aiyEpeYe4jS7Y6HiLzBUeNtaAArSDyqwlRYSONBKvNlrC8AKIU6X15iT
y7M+f9cRp0ZBrvSqhfzLH84LKm/4wnMlULaqC0t9ul3M7J2cVaOjuWz860QHjF0fWTucr2IH7bGn
dVNV7sUkoQZOJz5b57IEkAv21rqE598a1d9olBqWwGG0HDa9WQD9gvHaZUpH8n7L9oIdc7TZe8Qd
wnb3xaB+lMKvg8K2syJMtCDF8iD3yvn8/cr2VNv/TxnvcNEym1n/oPvaGqZLRY2z12wBbX/6/ptz
ORI8fvq/cGHXgscM2iLHtQoPrgxsraXU6DGOiRRtL7bBpa+eWjWXmTrXQbo3zSzl+nUbqPMCxMG8
z8y2wJOgFFr2uJG90AcecO+8+2vFdggRDaFswxgIq/sDQeJslabr2gkYAK6znwkOP5/2skBIDl4n
Ltt5RQ3vfywua/OhZEQ9lG6czCUr0z2sRf4iCbiVLAxiRZ6ZT3ItDGcetqg2KN8X8m1+2NT2vbI/
JRA/pa/7i+zxUSniTyQ9pP9QeV/VwoVnnW9tBuioRNT3QBdjfKesFIaz0Bxi6hJZgOzJ9zS7x4ga
CL3/i7Vrlf2zOHznplEmDwIhU5bdrmnKFrt2LQ3QfyKgQki4tvt9gQnhauyAUwvFCa7gNeEuwrFN
43d09CDtcCmvC2n0AmSLsBNM8+Xsfp64Osj7av73K5ALAxs8V04X9QMQNfZ6Jo2PR8WJr/I0RzCf
fN1sn8kqmodA+4OA4VeHWsNPWjXCXaKs5ss4UIeLqGpT0VTKM0DicTW6/1jc6/UOizugh2ph/bb+
FJiFZx4FIE48Si8OGITfkxPeumYACAW3eSohSpgRhsDmHcMqvEfLp39knQ9ZopkAZa999f5Tc0ZM
OwB6RsukRV7vU3CuAmS9NnYVJPF2isfqsMcHhlzj38dy0QGo28BjJaH/ntdgI9DF9/8sCdqeBJbC
xafSrSkcOPiWISZPJWcxlFjcSGz4p4pZDW/YR8jE85+AzvubcFXdhkC42mKMqWaVdgsm94WbVuHC
8c5yuxt0+htd3fhhthGf0A4/e208220waUTMZy9NE/QB4LLLGJfLgGWKP35PNpeBf+QT1kaNXpgP
YqoEQmODwLEGLPo+r3rZ/jjMCrVLuez+afUiAZgLiTdBaDWfkeuGrWWTTTnAv8HenlPYd6jVRT4M
o4YudBWpnSeZYBe1kTjm90t0U1CETwmW9uFxrT6stL1OWJ74TS6g+VvzBdBMGTW9z3uHqTz9weUu
a632rpK5utj/Jv8E7wGKh8FM8oxFZ5tJWvHZ9iMnKfdilF7oDb0iYme7HASyb8ndySJfbCiJrq9c
X+FOyBNjBy4pH3+7+crr22+4yrxlrBtBEXu8TZgfUYYZzbTpBZhoPDnrWdUUqHzOygnhMUCmFue/
vyTyhgcexImvVJ5v2VxoIeSkKJn0cHosGkY80Vlp3E7UqmEjj2b6Ohj1NPcRcGrWZDwzM2RCq9LW
HsO0VX6u85GBJaCVg42jcCMzQ05EAc1IqKymPD8Vk6ydvmfUp+GV0TMPisqGjQLGHzNwfgK46LVa
x4OMSoFSHi7DtnYNL1j5eyqnv/opdqYGa5mLxYlmtKI4+KD6uL7okenq1OZt8anORA0lXq4mFxwV
GYwjKCrkYY+RDG85JDckuRT6WxJ6O8X+qAU++dISknfZVcYkgIvfD37Ocq8upRhBO0Po745uObXL
SfHWjfSwF3TNxqWy+N/o8geWuqIT3qwwnBpYPjNlF9L2JR1VehZbijtgFMBPGNZjB6amJ2Endx5W
Yb+51i5YdhuaG1r1mGrv70LqDo4fY1xmLRoKTdXGJpzvmJc2cXfrfEFnzUhakSd5Hsh5kQ7kKiP3
EIT7kv7U0SUtxSaT15wUtMJgCGUOIlSe+Z1ejf0C3+/X/aMZ1A89RnRMsIHDqQEh/dQ9w9IZcLXY
DIjSLtDDHZNAlwCNHN2jdRiT8ddIrOmZdJRXrrAW1SZ2sKdJJn2DUzam6+ubvwgq0sxIrhtZXEz4
/B6X/LbogC0BHSntCYAddH9f5McfKJOupcisuTkejdG9tm0NdRZfibcW7I8BFV6SQRAoH7xSDLQV
HEAIec0Tsu0dn8kA+VVCaV8FlF2R95MZ27NsxMso7PKlyOQk05dqjA==
`pragma protect end_protected
