// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:32:03 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
i6QcNvcaEndfG5ZX5ZWo+Pz8wUP79liJa5hk1veabWqvYZdNBu+sm94g9r4lxOqg
bqJ5saPfGiB4FtSL5bqjBijjh6Zb9lASYby25IKbsT/iI80S97lU8h/RW6oZ4T+r
3ixe6bvLadVpJmy+nmHyL5LSOW6xRv7BQD+UiOT4Q8Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 58352)
wjTDuLeeZ0moL9PBzpiNS3Q5UbfyqfuKTwTYcumm1OU2P4Vv3YdnOek2XNsXpVTV
P5Unm0R26AJo4MO6E1zAgpdMIIRTzOGpbMI6fYfhhzcWPep3Z8OgqLFAvonTmA5V
WGKRdbOFSJmu+7SlXDKrkThTDQyFm4o2JMaf7kuiqZW5GDqEWHvdoZuegp6b+C7e
fMegpJaqgDHKn3N33pYrKD9dl/tcKfbtfOo2xu0YFoBt+kMOqTh+l0TKEN0dE+k4
/YJ5uIQO2M3doyUlsrZjSotqasuB5WDpABAQvRf83eIZuOLdbI+aPaXyRmqOqHdY
0lG4JPrLSjXiR1jOhcxMZtFcFPcW+Crci0MIklvmU7SEttnsYTAQGRAG7Lsn9Uw+
LB0eN4HCFgBabzfmrhvRGkiYo4lPnCMRBoP3GtdfYAIXaE7WUK0gJDwxqGnp2ujL
NYJktemNWv/yEROf/nQhXm90jw7T3RIcKKZyfIe69774C5B/hLOTLFBjxQVqFWVy
6ThUPhmOn2tbOF+Ih4g51pYag7LgX92ZXhOwTb4pZH5yjn4yrHwIi9Ltv/QQgv3V
YxLVXwx2/VxS3mp+QEJwl4uLEgktJjZbCHR94dIvLFlaqWh4gz/rM/EFB6+8+qo1
3sphQ62t1OwA3lLOpLcO6V0WoD001dYyWmaiZRkM2I5rBw2Uoc0+gWMPpnDIYmUF
CUK5g7J27l+4NMni1R3TIZr8EmB5fKYtILIpAiF0dtQEcmWqMSflNk41PWEx82iz
jo/PsOBtLwZslmnoAk1mqayPoEVLvV8i0cSCcq4mhWtCaLytvAvWJ70+9XwfYoHn
kBMLOaQyq+Sy5RixGSd8ZjonPxI4qOQ4ozCH13Epi/Rdz0To3mpOMF0EVRmGN996
JjTykcFRfxKn1OlUIxtl0XFD6xfSFZ57qAZMeHmwZ+G4cGf96bHzZmaqfw/+JENX
Tw6v0Tr4YdJOoeyHhbG+0gwQy2Q/zifI3PEDhoiCrcFTxNr7RkLIeCHMLf6dwULQ
gHv/gzGuVwx9KEmNq5OCxrgHF1JW7b8SGLHAt6zRzmyvXDTrxugni/BheAYPVeVA
I6FxL75ymb0sI29cVSx7do8N1NNDIM8hORwYZDHsidyUzoFKVf6V3WgB2UFkEXhv
g4QqVM4MLvwC3oE4MBL30r5xYBt8a8PQm6Ol1QbgoSoTV9zpSh8nM3ewqObLdoJj
BEfIUAvJIks3yWk0PwEcLZ+xgAAdDOMZqotqakumKVB4ZQjYZ1uzQ4T/pfsVu6fZ
MGx8P83WOP77MN0oi+rAsqoal4VvilzuF9lfBWoXeRGP+XkYyCTEkTTbs2ZHMuX5
fXYM3hQiVsAxW952VqK7V6QFk8gFEzqNN1kTg8chdZ6eNtXJKpnfyY8lQFhO8SEm
RPGwhY7T/xkhyWc7bR7f/DNzjq4kfqSzO/aT2PdU/dABH/Giu3SsdNAENFbIwu1j
X7H7IHz+CmvQevgzvbZd9GDzbfCq8soLv1rUyb43jsN8572LZrL8DRdaOE0u83vJ
BwUchv4NuKUP+c6zP/1CMyDNrV5pYE3vD6VxV1BC/LFW7PvAWnHmQIXiVeNQI0s1
RGPohngnRFT9vJ248OvFSe6/mGUuLvLD8JxQWMLgbM9bziaOCYuLnEkWCcsFJggt
CTNDZe54wvs8J1vZ/joLEWhcrBfWEGndAkIAj4L+uzXRx5SZjNGV6XHfSy1yrhcm
nnRbRLpRhGgwfc7a2icvx+NoG92lqH66uiyHwj3xnRv7hgkwFuxIZgMWcGhQECXC
tAJYbcdi8KbRbQ71PBocisrtm5Dju6x2Zi4pjAh1QudzlzNkjAwHhORLYxnU53kq
t6Nm1fvyv4LBXEXjnUM6EhmHPSCVxfpPbDrPbZ0ITDfgzMNWRAanV0w3HEHjC87k
1D4f/43gKkEa9j53MHXucEfSJVp8jm/aBQqjPKp8KFMI/ZuKvL2HtAylhv+M9NrC
FzBSoveHEI4795j1mavmqG4qRPRgvSkMSIls8RLBLG338HbcEstRkLgWDL0fNaC4
KYzCW/IabUp1/LkbDwnfpASn9B6G8u8+caUDphUQSaPx1M9xAJHHaq2Pv5T3YBxJ
065OzADHnfOJvw+pR8KcUEGv4AznJInjtikzrgcQFyGJh1qhXIPo26KWtkOxp/CH
R9k47IGQ6tlfGTo51376e0puaYZVOR7DDc+C9DWGf109IngR5uOSFkNG4nb7dZo4
r+ttcRLc4CfLwcCYiFxGRo5B7qRCuFvOAwwduTpcBoshMNc0X52eAiRhElascGH2
kmdugm722CYvNTNGf0bTUNpoQRqA24mKYmmtr6ZOJj23gRSoM+byxI20uT3DRUmX
z/po2tYbSShNMWM5hFFiMNM+MIIA48Fhksv3PuWCv2rTm70+l3MK8n4TRMWAos3p
O2reCXcWrbBcOpoXwWkN0oz93GNAHfl7A5V2MdstzgzmDBXKVLH2vFCiYWm8H3jp
Y9+MfrhMneOvdddPHNFJtZLC1GH51qGPmY0oPYZr0Z0UcVgzYm+9DT1k8v99Op/a
eNDwCkgpZQiA6N8c3ujam40iiRkHpei4mG8LIzfPelkAj4QPhKDolK9XjIrTMrUA
WH8nXRMgf8KiCzrz41gswiGzqQv6Ek0qxS9ECrCQKxy2bGKk5pz3k2v9l26saZbJ
1BSFaSbarV4i6BUV04f13cZ6DMnIdLCpxSbS9R1o4aWXbQLo0tkf6Iw34WJZCFvl
HKlyEbVkiJZ49OSYY6YTrRYIqK+e8A6dP7J9NbgfeOZyn1EoV/7JW3TwIp+ECVo5
jr2PnMTLxzpica08Bne6U03w6mcOjLtj5cOWsSyQg/irckk93f8kseGRQ07ddfT4
DNNuz5UrArmaalHMii8EL2xayFqFArniNlPbPegVegoaMULvIXm7+8t9YPQCGnhs
c0RwxsBI/F0mFADCkl4eGds5IfXKnTywjN4bLzViuU04kw/A3JYvRCPevgrKx7hl
KOlaePMQw8Gq0nLAAbzm+u4Qqf3VUfhAD80bD0jB4r/6volsNjvhollZBzKaF67j
7w//avqmk1GSXHo8kcqyhGHZwEj6I4K/WerAH2GwPBJj81ct3+tuHijyk24sc6hY
+RT7+DM2s0bmj0TYcvMJ2DrYsxjhq8A/MELSHRwQtycX3AT7w8iJLu0F88xh9ACO
3a6jhQd0EL4qgdV/BLfHZMqh5I6umiHHpb7plHwGUx4wghwTR/9h5MmzDkOU8aII
lYxNTKoyKEIbCRZHzXAwKWQRZhHBuzTR5rJfK9IX/+dmetS3da7WwcSeBzHC9YtS
EtUzNGmCqlISB349kFZT8BSWFyN4wxKF7OP1LlU8KZ9VJm0kTgcOmZvYC+BKxKxC
WdAir7j8V3MT3V6PpY26IPF4irpL6ZFQiihGQ+GmRxuhg0/92VV7yKE1cpoMQYqI
XHdvSTKKthlaDOzblydcHlboIzKLbFedj2vUh/x00e+TMjnMkYpg0Tn8tgdB+0qt
g+YlR9bQ3lxYFMAETjMQks3r6Hj2dnI3H+skXVqFhDnKgxNGJFizlzmTW010GNmb
LwlVXWzcSULyJ/GppiTqvgDUhrHCY7OZFXWBbuB1ay0ZPkzRe90MyyDNUa/rIJO3
JLB5hCVhjEsVzIeaDt0EBvx2vKsxKtfaacMWI/JPDOmwG9tGepV4otnJS2a+mbGT
ktOe7txwc/dn4yQtTzgk8he4zdfZt2zrqNliy++NzgU0Ydwq+n/m/VZjRbWTNzfO
V/5yinY4qWce5HXtOtg93LjfikM8AyRSf+h5ipTL9++ohOmpMfj12nKUDVHpPF8b
lUc8o73PP8l6P07TvOocOVqgQDf++5JAEA27I1Yysfsu90LfzBVkkis8Co5BeudE
Cmzan9XcKfuOaDUPJBkXtuzm3R9273kvGRjevo7eTLyzQVANvVYSlAx3uzZcaS4b
e8rvmsX+dxWuiTI6T5t3Gd1M+m7YJybpn6k3MrL6ZXQHOrj3sR6jAeYaS7hQSyIP
s8Lbtr+nQrN72ohNcoCbyQ0CX0sW7j5WZ+YidPbCoIMpmLPPq2vjHbJ5WPBPPkG7
ANA8xavzlARN+UuxuW3OnKw9TsPUdYO3nuzDRUW3zSCeITeplm33/g7kSUdY/pW5
zVftX/T2b/jcCeovW52lOiZaGt0s0bwK0OyRwTuT6c1Rx4Xjmw8CcqxQrU0jPLwH
Mb9Ip7aO1Kn2gGc5mHQ+Dux3tQx+JRMOuX/0BAwnVloCi7piWchzfW2JZuqSvP+W
EiPy7kzNWnhuf9nNUVFAIq51g+Ag253WKcoK1zwTGfUM7a3r40sE5RJrpI1rF0ht
9ebxQLvZU4Xj2Ri6SIw7w/CHya/zMabaiaSYHBY2AxeBSeMnOnxeT0+dJmwhfjvu
T5WRhhZmPv3rJv0T9ipD3/K9yAn4+sNx3esbAH8o597OTgtX6CQ+Kyp/CqjCrEpK
A4jcxBZOq63FffWr0HTrQDjtSi8mxCr1gjI/kc63EXAGo12JyXbbAeeUxF6ybvxF
PVsmc3sG4I8dMAHhnZMIpFeI2a8BwdwZw/0BE2nqxCDmSGdvwqq5B+z2EG2+nZQg
DFXBMNu6bZxtov9jllmEoSrVMJNLEcQYImL6UiZWPMjBinRPHZEpOxVeFoAoNgEE
iwt2zMSG/VmHnUePXQQAKKGPXn6J8N8CodHtVJk7Wk4Nv9ystbEpeabP1C5RwUFO
TrecChirOWCdlTX8dJofXwJsN2UfjoKFCyO3H6aZZHgx8Uo72oO8Y6dWDNE4vGJj
8VBnV6TRZasseMBuQTDu/AIkGxcbhciweOgCitZEmkOCW9N9Qc2FKjxIA0n5b/UB
8f3JatrjAI/Ni8FpT9aILlIF+YRp2+V30YgZYmGKiSeJutFIHsNm6Ejkam08L9xb
oYcmjUcXvU7J34bYWVEn56Yn3ewjnr5/cx9Kw/5DT3sURrH2kdo7Y12l1sV7zOvp
gVhsy1nNYeSzOmwBfXPE8g5/Zs3M8fEfnTQbnitVcYWxS7OCb1PZ8Sda4R4z+OkT
5QIrdG8Im6VS2/xpt0LwozP0v84jszn7ZY8V26Ewm2YCO3HzdfO9gp2T1xBf8EY8
p7KkPLv9k69tkKMxHyRAI5Z48Svlo33s6oz4FQMtV1ghuEQOiRdJY4gIQZQvqKRy
yTiWkuLJ6VbOFNOihYvesEotVn7BXSAj8niyUboStZqZwSCeGryHlH9B8A3tT5wG
PF2WJCl/uC4oJVYrwnoYqgbd0jLJI5B4lmc0PWjfCRQRps2C3JrLO2FACf/oWrJh
uiEiIiK8ZQeryBlf6bTbuTv1S/ew6Sc/rJY0reiqbg+xPoxhkLCmKC6+mF14V0HZ
TuZTymQyEnipuJpOuuhWOm6p1+Sj/f4M10Ady9XCaVjtFe8EmdT0/iD8en4huFqu
b0Zh2ZpYIzoJ2gkQYQxWH0gWbZNactfBUA4RlO38Ot4cQREMC3i4KVklvnIwAD4Y
6D3kQr3HW7iL+ggsxOmo+XthsdFNX7/zPQ43NdPQU85xItCTHx5jP4FW50GKQ92m
jhHIEQqdMzlBhmtHBXtzdhDXO8ajTjSVfpZar/kcKUQy5TGnnRGu8RF86odW/Q6M
rsvTLa7OBRkiXxgx5OLTiowSUPjhubP0J0sovawBpeK/936857gCKK7WZsMYmTOz
+BO9bnlOcxVPRYP1Y2lddMqdinlRuYrC3hWLYlWONevYbMYnnYMOWGR/Fg0oQXVl
+f9d62KAoHMzbSrK7mE9z3Pl/owwpjZIaaHBQrE30pxAl/JxgV4kzUEOZhahNsR2
utwGfiB6oENdd5OnzAfjdRd8j1itXMuzisVe7qQig9RrfUa2KYHOoGCDgMPoObkn
SJaTaXRa/QC3NCbPNM/ZXseUFyL5DZnW8RDzM38/LQr7kS+Nba3172ldP4YjE3tW
lcM0/1hnsIOk027Q/OcZUJsGlkZWo3dRbiRV64UYRGUP2uyxfFS2VCfz8bR626hS
N/niPSUpVyPIXlmWpvTM3wGtiliNddmcJpRo1c/kSdb39sqEDcYN5D5+hkqZ48Pv
K/v/2T9CKAkpPpSxCNF929iWJChMR2pucT2FVogXVM9gegkUtvf5PR5rSV61RLuL
XfLZT4lIN2AnQ0cmZ3rMEKfinV6Sr2qrn1uLSAt9YkZpz8NcW/iX44vUU1W/iAXm
22/KcHkWTd/8vN1Ob4SK6zkZLGyMwTLCte1T+ERwsiWrf5H542MgKSCAFM2UiyrD
EujLFcFXrPO/4PzH8j9Nlfea1ioP0V43qMVTx/4xERWk0lfPEe6HPtzVIRl+YKyz
hWvfmvxeEeHO0ARYDw8MImFU0kGf03i43ep3dLt0qebuzRuE9ayOInECt7GcEY/I
XwhcyIhtRjfldM13FNC7SNY9tXmC7n0z6V3fVxE/vnHgaSnX0VzGjlvC9EsLBuc1
0mRVmLNV0qHrqKa1K+TVUrlAf6fKkV6sL9EBSdAfEgu9QZC9NusokFV29h3O2ETM
bkPliAYaJIjgxEFs3BnI63Sw3vMG4N33Twh1rS1rD25gK7LsRnTHfSKzds0GZ9ra
8xcB8/CUIh1Rr4AbopWR/MAZ4zGuHGYu2eX7pHVuZgCE5j9rz4HYq3/JY1FRK0RH
LLkrAfpwx3RjRHfz3UXi12QfXPpyB/9h93s+e8x5fAJ3Xz/2PuobFhFM0izQaI5s
mizcVeNd7M1QLLwkEh+qTwuAV+bTR8Xs26RQGXEqsXEn4BTziRNqr0QrDax6cb2N
KaIGfaQh62VcvVs8EAWZTKD3563T4rrwHgHeYVujePYH+QJRCuyI/qw/Er2NIdUE
csvQ93C9YIKb//k+6ULyv/+11qWEmhKbSSO3UpbK7UpDyHxbGgxgBaysotGw5FGG
1JDf2/fX7UHkhGMjJarFc+LHJSuwigLl1ZSAuU69ILiqfiWGnhDoq23SJord6H6m
qlradN6iYGSdt1p0lrp7ZcLMed1xsFtwPGV6DIiTJy+S1Kj7cDdN7e0ZRwNY8EmE
ADSEcJYhp9Vyk/Uoc/JSBd9jfT8kUzHO4jdTenFdzqyAAxShLl+LxjnBGIHPiW4m
c4AjeDIMpGYbm9BNhU8DTcoRKNxvhrseAPDkJceWlPEkn2EGQNC+OY1yfzDI8X+z
lJWfnFARc2ijmm6hWwJ0Ti7FET+XUHE0CQ1nOhDDQ+gVnQV/ctvZCopX2A5vDFQz
7A+Iog5eZR6WfI7waqTga9cXNObTgtnVOBeNdOtLrVCY/wRotzdWvfMjVfyE1EEm
B/A64o6ooCHE9tNLNYpS7Tllsund/g6PKZBfG73wVqQFbto5KUbkv5zv45u6Ospb
phC81TUwSkkr/GypTCSl+a2M2wpghhlQEoSIxJb1cs37/V6cpH0cNCSEVeLBKXch
+u38iuS/czwXTZEQDkYMDaX8gNG/r8RZDb16x7zPtxPovd0fBxDmsmxu3CSY10sQ
rP0Qz/HdlskqorkDkW/Owb1jftcM4hWDlM+CLLobCHkIC36DCoSc9jt1XM9KEx5i
q1674ZQ3LmYKgqbwrzDm/NSfpLc2lofWtsKa9K7w+mfayCf+Y4+zCc43R2jiN0H3
ml/fxO5OPKU1N37WPF7jJgifOUZRoI1nZ8ehD2HNZGVHM5PODQo6wrObyqsCTSFl
t5JaK7eBr3nhyb9C+lY6MLtfoRoBcmuTUGPcAo5s/E8mSzkFyvEafHUHvIpcRtoE
RWpdhbqkhCATDWwD9leDrJvaIddnVcUUL2leh9msXdjBhGlyMt7pT85EDj+IFaeB
MNOBYEU30YbMthQtfm3ssnPQIGw7zrsgSSVG7RLFjKD0kQZX6/LonZoOa6nO0+o0
z58Z/ht668W+ln1DVSEdhAF3Qu4jUWksqqYxO++ZJzS9psM6g9CtUJjCorXaTnrn
Tko8tC2Esi8h6BEuEofJbYfCBWpyqmns5n6GSeMmcu0B2nemZG1mrsJDRBhoQcxN
MxGBVFerJ7wu6M6iqhxyIZwk0F5H/5O42suDMxlo8JXChyTpZZ46udj38mNP3szi
YytWF/hdflIBnRR0joHFTA70nghGbBLyLg4Aj7rW5TSn5sAfuPj+XfV4hCnUBsLt
nwxs40JpDVkhnHYhPkzf/6l+2yCRK4yojVKDu5eUlqnU1369N+yHpkaNrw27TQeA
6HYQSprDmF3WaWFL7ojABcdVHTk/PYuZAjdWkG6TSBOzz+BjoOfdyZMENTHWcSTB
xUi5hs1mmZgMHPUPnF9xIFr0HU+W+KVNrVb6tpOO2lOPqjO6NRN57/M9i0bkLMAc
91B8DycF7utN1JQRy7bewsPKQ1LNLrorQ2/quk0JZYOrWnw7OkRVdQ2YtO/HSiUo
i8LPn5JsPP3b1kyXnmS9fL1mhdm2sQEdQwNjXb+ImVIDqb9VIpk0z/RHb5U2h1H9
pjGIwD7ZfN3F98+iwlY0aNd5/TQ9LqmtO9IqQXFl9QRu1KgNm4iE5AKSYvowa8N6
RoBVd8tWB3S6JAyLACjiNtBXwXLERQ3QGJkZx86LVGzTeAplZkSTiQ7IlpIelQew
TQPif9uehSROvXQcLQdVPIqa9L4CbrsqFyjXNBsbqfYkyl+/Al8h2UHRJ8PZxFRm
cDn7aRpXSzU20RlK5/f5W2I3BgllT//5S78RQSXRykGjLpKWxldUutK3gM5JyAx1
j4rZFwOOINbI8Xw80q4q28iC6sPWpFF75YW65ZI0FJlWHA2ACmObQINQHvrDqi06
+cRkthljQ4PB7mYavu9JoiSaUEvIeIYx2CchSZRkOhQF02cHz/6H1Z5FZSnj/tBV
7S2gcsLrh1gNKJIr9ZEszGTvJJEBwp6iSa2Tfi+n0z4byeYP7o8PlrhnkDmX2t3U
AwO6bxIaywYE5gTWXOJMd2QW3Lg/fJHQRMrcFRvoC4jBqYoHvNZGTW3eY/3p+Hot
oTtkA5lSq6VEsBxaTbstsrnTMUd8667LNw2T96VqllHzErACcg9eEfC7MSamZbcU
Wf+fz7Kh9jSfe7yqLLRClMqt07EbScD1DDyhK06xSZY+TtJErzrMGt7Z3D4jU1gB
weU4X9YWUeCx7HC2gq0ndw4ZcgRqmhQyy6cv9+mo/Pu68KerEPd7vW2onC2/JMkr
+oebK3XgoYLqRv0IHaZnMUL/VqExJ+O+U24OWrSS7tr6rteO4oXK+jph344Jl8NX
rVhhyXyvOuPhqsW1rIp/9vJNuaLgUzN7+ExVTtLq3uuiiFhbfFEr5578FDExzlJJ
uiGGYjMAzaRc2v/9CrSpkZJ2SNj0/8ZfbW7p2+vMDmumaa9O2LxViHMRwiuj6oUh
B0nrQyELyufU0dv3k/nPyJEpN9NPdNcQz+TU3oO84tXMrS5qGkF/xbZewKfkMhL+
3ShjCH6GO/Hp1Ry7Gmp44LX92bmzR/s0IQhfg+T8SqOQGgYtDIixT4gQlmlRTdV+
iC3spQphJdWDwH+NH58cwLbvtyxkPwx6xcEzpQ2HslG7Op+FbfyzKczks6Hh/Ycs
fBAtwZZJJgMIQ6dlHzxGoLjpWScXSRdDTNETnx0mZN7ZlLy8HkLJjQjphKu1biRh
196X9eYXEzU/7M9mAvlmyvuX1cBjkqXrUvEOdcmBIuhs9RtittHF9CQflHDsuXpi
dPIf3xGpCipXUIrdLhYigd6wima+8L0AAlYqlJzmk4L68yUF6497WGpFQZB6HBVq
pcId3xzJzj1pdFGyjp7l4cf58RwaC8sq8U1Egkd4pH5GvVgUy+kXpTkHJQD/jRpr
g3oB5PtoqUAdc3C8SrX9fMnR5pACV2dLJPcnRHCOhEjbv/QLjegYSYY47G9xGX+F
0JWW9TIv6e46/ObvbS4hX1U6Sr5j5tS8S/sxbMJa3JSo9cm7hr1NDbj/EQpw5Iuu
WNBXR/EDI20+k2DKCTJPunk8cvSdv7Gz1J/Onka/5Np/GlyI1jzBS1LyDNS1zSf1
ZySZJvKpq1AY4MP8URgt123zbbd/n1DvPAzd6go8bjV+c0XWjPmF71DvUJIv3cuH
ZgUrkS2GmEO2zHOfbTQA8txjFeCiJSZyOg6L5GDuoFcneU+mvq5O4zFrz1QJp5+h
14r+a96arR5zU/11/a8LvtPT0VWgmYdg3l/1Q0yHL92nlg1JXPqORzGh5/EuVvRJ
QInoPjGUQ7zgJKUDOflQxXLcCD7wegJ/X8M+bOWyZ08qpUAC0ttOxJ+xRmDkMLdI
+6T7eOMVIRx/NwU5kPVK7uRzg2cCP6HWb9VPcOg/g41bjdntWbFXWp7okoQisaY2
akeCmW37ul17/NGitps6fSJlLNS9BsDPR5QYq+HLn6MXjYL5WVdI5wHCzPMqej+J
OheMzwxHPuGzUtZWBcGSVaCrntNuFUCiOGTNM7vCcRDSXhxCA8Ag/dRKK5W9fUKy
dv/eJ8W7bEzRcprpiaphae3AYCe29T6u8v+P5RjxJW+20mSX0OU4EAdlLUnoFT0Z
UuC18OPSDXR2/xpwiLSgm8a7vscaiuaPqNxst0cm/zVniZZ8oZLo5Cbzy5ECkCgi
nTdgmDwHAvhJfpkVHRtK3kJhIwPX+vCH3HVsmV/gFqovAxeMKTp8e5HCdOrc/m58
U5GGuiBzE161dvayg7YLIIVknh/RCah65hxUNAKwtV9HXA0ewpjZu69aNcQP9a5+
KNQ8NXArdwNYIMvXVYk5YRGrJ0SkqzHiYcy/toB8WeFnE12UzJnP/Dttvbjk6Vij
hMBQWhndJxXWCTBp5toBAV9xfC1YAre0tibupFeJxtcb6QFyjS69WxAsemI+LCz5
YJOXUuFrJfknRXXX8LifsgqvL3r01NmB+WBvPh1fJ2J+3gCq1xP/IQYHmiUHjjz9
ej/45SIYzE/pPHi0yEkLvIb9hqwcX82NEpQ3B899UAo0J/JAXkhYAOhgisJTXbN0
dr8eiCheUMXnKp65C2HdzYLhlK+odVyqJTMo3CmrZqWKUejQhMUrCEHnD6xwvc0Q
QHGMxjsdXHD2NJvgbqL7DFtNSwFZnTXjjJG0tBkS4F+RnwzhvKTG/zr9mPTF5dG/
Veocby2oq7Y937zH1nyZ8I1Q3IeAS5VUw09VL1j4eJX94EwT27Mab8b6KYwnpncI
aIl/mvlhn/N9krRMnJqmMK7ieEFR/fMv34zLXrOazik41ecVbZavzuzhHEQHszWA
fUXuMtVaKDWfH0QNOhYwoXRI3vBYivTSAC4AozaFppWlS9HZzk0CvDrO0vaTwH/B
W8u1sMYLXYFnmasOpFMrTgeDqnE5rG7ze0n3+ybvS6HdS57Tu9h6GfKSc4v5TXY1
OtKOvl1lCCVXbufQm3RZkRuHqwlF0yspH0ezrGg+MrEYsKn5PQIZ7VsEWc8b0d8H
UHyJq9Kz1KibjcWXmr7BuFMtkMIpgya8U3HVuL9U3vrlyNVxEBtoFtoGLcP27vnP
PGrQNjj1ydmcHzZi1I5kNgzm0iSqJ77PEZqTOWKqeHlH//Ba9ikBK/578kfAtaaj
gHmI+o01Om4WJIabjS1X8j4MDv6vd/tp4a/gyjQO+SYKrGTy7eMD6ZRmrlwwG1sC
zczzYz0bTSjQDcGhW7Sv2qzb7uDJRVXY1UAlMkI5GwwJ7/oM0Z+69meaKFkedtKy
RE1bCqhp1xYAosMoaHgQ+0jaLpa8215iVt4F3dAULwVQh8zQZVFact2Z8R1wKJI1
ZnfuwAHrwDJss9K2zULCQEou7nkXDR1sdtNLbe0WadrUtnztnE4SgGIpkM4BBy1e
dBwbG1n9c7a+JUEQRsJ7HD+2GAl2Rd75Gq+S3USFSb5Nqli7MlpbYOmZqLw2Xn+v
n1Mrh1lLoDDkLz0EipOx3B1/BweecGsim0Ivu/5XNx61sc3YMlrjOiUkUJLdJwK4
+tV7WnAEgFIOamelRipRiTpuIHtsr0Xwj4NEbsTOgUCnSOGWKD8tMR407WqDMYP7
vdi+8YBioCG9CDg6SUo151SQ6WdeFzmE/5zcyQXDJEMhDxay0JkSbz5CiUnTBRme
rWFE8LJw1QcSvBm5pDA6LA+p6RnuIAD1X3kAihU+oMkKnHEr/NOaV95IACB+VgMp
zRG1rxK9IijJRPhywoK5TIf8JABwZQLQ6W5FPaqZyN1AeMp80ljbpTFH8uPA1xXt
IcHYCfginUYIFAxO/nB9FGi+S+c5ESlMQWUHtM70hpuD6HzSPo1s1RhcMzQijyBU
CZNvb0zvrpDwW66R6CINmaQjhNYw0dMKUplyHfZZ3ctjvCmzX5QP0kAjmxUPemdC
5pZg15/w8GHU+Jz/Yf7MBBQVzaLgEvarCfP7hFbx49lbfZe0iVjjoGaJuNfpSpNk
HKy9qCxtSxTiNTr65dz7UsGxUkuJu4otH/8SXlcxt5JkIBPFy36kQUYKmdFd012k
6W39vE72PUKbbgx0D4AfC7HgstxI6ty7CUQkVDxly5Bv+i0mDgglvUIWPEQVYNN4
Fb+GbKzyXsJDJIPoV8E5uB9ztHRlSZrV09ehs38kprfw0KdPVA6w1HpfOr4WGaB9
FFPELbwN55AWmCd10MkBZ8BR/YeRC895XVYVlUFsZqRXY/zEGY4lxUBceNmzE5EC
qGWp/s9Bs7qFWxiuTeItJaLl0Qwv48bf+a2QwistajHIV+mzmQ2lb6Nva5+SEUdz
Ut3oHTOHoI/kG7kWTRoiqHcuP3QPreeol97S/VMNvKFITZ6dqRf+UIwOjSWl+g+W
mjxXSRLxAzcos34qspJENMsBXf1HGVGV6kduK/G1HSs3auu0PCmLF/1avUWRjVJD
XO9IAlpOVn1sDn4wVLWiA85eFQf2oG2or9m0HBSoju2Xq+SPhv/q1LMg6JpWT6VN
jfhAS/cGy9kpDRzXrC4FTfSER0GzIV5MsRYqFNLaoO9DC4qfXUqq90up98uNz+IE
U/xqBH/RPZfc3EX/Hkgpa8VEXbN6pl5emMigL+Jl/GbdsgI5g+N+NkOchJgoRn/9
m62dPA01b471UJpWmyTWhiwXH2WNGK+h+ZdtpTBHQSsIW6VSyWStT7Rvsw45tZHZ
TGUXB0vpLSjGrlEEi/JGo9fhRx2YtW/CvMwhBGwsIvOlo/hykBJ6yyHBntXiRO1/
VXbrS/C1kaX1L0EWtx4hdA+MtRSmvVwESkYvQME5Tlplm1LCOvJ+o9AnB2SIUZIA
EmaRzno57fHfdB9wKjZyL2E7O9qwzvi9Nw4W8AJHbai/4JbUUoIpE7VsN8/TryNs
w2RYCKt8zRhWbDreayn0Ppbv3AzS5JVqXEMW7AgyH7Wn8l+LWhwIywINjmqLPu1H
Ocf/PmTQlN++b1lep/P8gIsukI8FCQDpfHeWVNb6Zffpmj5+Wlsnqj9nUDSREutH
b8RWCZnRuCxxVM/JMRTIuSLtnCQ8BrfC2PWcoezH2kBtZj9PmmoOBg9o3Il49aUR
bN/NHseBg1iEc5M14CG89GWyXyRIEforgUspZHRsSgR2kktW+YytDvNv3VPfdqAu
chbDXkq6IFnoow+LUqp1Wm5a5yJegLplWNmTgPjm45ZYJsG/kFXY8dE9TTl3mlBw
9uMhTG81AlRVMlGRKjK/oijLYq9UkpB/d6+MQIePTnsNSC5F5SekJjJ7ZfyUFT5u
z69I2J6y8ntU9Z++svKgFscr0U706mFztZmgOSVrrd0AppuN04rLvnj4JvGLbT4C
GZUJuampUq0Im81c4/WxxE4p/+/+bHTAixxNVp7CYkGARaFMUrQXEErakZEALhny
NUXLNK5rWzGmkCgvjalnmOqsBmgogkYOls7SfRhmeHxZrTa/B6yV4dJaMV8DYAYp
aiwHKRc8al7UWB1cOMmcapCC10IQb/TphGwq+m6YsehF80ou/WDDil5nlPkOCeik
gk8oGHmXjAu1R/Yp6FzCyZmTBbtv7StTPt0JcqtbKC06tCqMuQ2NhqpXVwABEbRi
9l9EMfK2+SubdZhvQxzAwem+HyCM2iiJQcGxqQj5C5f3+jsxfOb6armcJ5m0nz6T
EUCXdiOy2OnQaGkmS/sWE+hAMfgQ2CYmNW7kqOt/mhLAM/JbB6AQc1ecqUJee6ev
28YyvX8pWTeRRqlaib/UC8KsgTGEIyYL8Jp48v8RqyWAB0qlstXB5QhPOL75Obd9
CYmrv2u/eIozPFwlCnOgAD2qJJdmjcPhPGxL04WfnpFarNo17rG78AeOw8AceIaL
TG4iiS5nmHKfepT6/rS/J/W3gMhmlRAAtd5QhqPwkqIvSrBVGRzCXG4ypdT1R0a2
vQeNpBC9/qPf1fN3MADk35rVqMwrGATgYTZ7WtrwvONJodq8qJdyElKdHmphKGKc
NXPfse/Fv5YB2jsOKC8wZQ+4g7iHYPGxlbWG/HVdvkx6IBRQ5jBUWL/ID4wUvFZy
gyHYNnW0SqX+Vsw1Y4nec29tNkQZUansYteBoujLwUO7mbS/XFSz28C3cvJbdzKU
fS+RM6hG4ZXDpwl09KvGNYKaYH6IotL2W39BrbbjNUaHPc+QNdNNBkaxlYlLL0w3
ABB9sJj+ao+1y6yEqDuVTU87zcEaXYTiLK64GfbOTQlDFCiBQfDeKTHNxmDMMshK
qu1XnNPzmWrQrTfnb9oj+VJJGBfSHLgOWCe7KZWGAgEauYO3CKjoPdhhhaMyJk3l
Q8e0Q4sYosMj5P4QM7Ig4hujxr7+uXnp3CB4HC0EMPMHedPArBB5Faznxy4Jqthb
adP/hrvVRS/OVeXcmeiR4fX1t9ytLpVT9V3ROERY2mta8ypc0nz/QcUpv/4omBwu
NVOFhfo9H9iwmylCqLIrqKQOicLbUMpw1dEpwETVYEkw1sDSI1c5FDxPdlpYJYfT
ZiCPnB+h4AZhrXFIbW7MmUpi+KSOZTjcSDAMsmCVuhqHDXTAoploRgYfuC1Ja88H
QTXLLrina/x4zwFpoWljBKeiOHgaLuQiQG716z+kUDS7TFcTC84ckZnobDeIZhzd
aC8G+l+1krkUJ2mhJPVkR/bf2cmO/y1k8adMPhA8i4W0fE4yscyZx1WHTOqnWNlh
MnH/OYtXtAFIXcTlyWFwn5gTzjhvBWVXCWAqOYcXo5SOkxMIuW8OS8n0z2WTLpUP
YR85h/Jbybm21sXgOgD1CQX/aIVuWd653FAP3mN1dVn0x73J1eDiy9GMSRd79dch
xblt3ihzfqdOiFSci1KzTQxfHtLfcKde9Gwwu2fhy7o8zAM4UlEpqMmZMdAnfG9J
nIyE7s/QXYpVo3fD4hROin+ict5Z3VdCfYBfktrqMydjFeayZTBsreDryakyvKDl
cApQjADd11NBeOD7ZMDWj2cRiEU7w3qDZptIlg9Nq0wFHQBPERX1s+UBdKRfkT95
NhAEL0Af64WmNpAVR9wA1gzAaF6A3qugoN50WAiq/tFxsPQ9THTuWEgLZHF7vpya
bPn5y9dDLzAxnMibQPat+xXsWiHDmrjZfMRpoC5VpmySZRNB1Ct5lFiqX02RF7/K
q8vJC0U+NcynJ3k0K9CKqqsf+kZSW/dIvlYbwGq8cXSDgDelLNkZGQxTnvPks46J
x1eAkl3fuk7V+x5WHs0SQR9VXxIVgHeCdH91bx4TF0b1qB/hW3cfTfI6mbB0JXNB
U6A0SebequZO5YFRF824PO/vRJ57UBpQR7Y4vSjJt9OLTcfRvvYe6rD0XY0B5wVg
SojqJR+k8yZzb2xwBt/uyyF4z+XZ3GPlNcM7iQZ+jOwSb5SVEvCLerIfd94XhL7F
qtW7KnS06wAg5P1kqI3Xy6pqxfByzXfVWa7kqqxobCyYVTUlCdHFDiDPW5lb5uSD
Cq6Es4dARDssuEkH2h90gxdcfeJiDHLx4ZgiUVKiqLWwvNqy/7k3BRFhKJWmOZk3
eBEs8BJtZ+qrmPY3zBbUjje0fQ+FNrGdGSMNwvEM7maR7XpV1P0U0vRwUaP2mJGu
zdeofGnYzvupEEjCYL8H9VIkdOI4IZ8gfuJgSo6FhyIHpeFLF7ns5xhDhoY83SC0
jbH7z9XnDL1JdDAb6aGwZreE9cN4wgKbcidB8bMOnhqKkfXbACdEQSOxCKFsX9I7
MEcj0XP2GRDL6Vk4QJHpzEHrknZ7Zwxy9S1Lsi4sYIfkNcslJPGzKA9cuEVZ6U7Z
NmSana3TQDMj7mVi6Wvka3CZSYoLTiiAeVSq7cI01YM1ZuGdeN+4LoZvuGk5HEm7
3cyUfphI+1togsflXQbCraGWoabbRzS+E0qPMKKoykmCEnfdmNq/Bhyosad4f+8r
9twyLya7fux3+vALZxFbv/IFXYfHLcP6Vfhx3Kzy8FdH+F0o4EPM8Z9hPfOdJt2s
ndP5WPQui7b9Hya6HXAP/FM4PbJcI3FnV2eny3O/JpVLCMInpoSFbhnhtHkv6Q1U
+qUj6VoB9wKjRctJiKBfT4ZYkPFTTGDVZ1zsZrPwGvhYluR0IOtchS2XetBPHTKR
LpSZW1/hXXFZqxYW0Q6jHxcEoIzJBUBJ//ndV1kzZvSAEuBBIv0iWajIpVCX7l9u
s6A2ECUggSbZ8CniCVGmxlw9zwNataF24sAa3/RurISeRSJxNZjEcKgmdRFfI5QB
dSFKnv8wdB8waKehub3+aKmPalW4uxSGeXU/XZC1uPavN5BFDDvn07qcxfNbPyVy
jIrMAmbshCa3mdUvakZVRP7yPJkHJtMMRz2V2j0DaWTirKfvbmjET9FMwHTW/j0O
BAZlQBno/yxLeUBt8w1QGvqDYk3oHayKdnmxMLbLs+52xkqCDWfPL+aYwdR177Bl
K3+syQQ5459GJC53EciBlQKcZBEK/+qIIfC/5g/4ZrR7tPC+OgjRG3nVuhh8u2ZJ
rf1Z5fF4bdwMAXy5QKfOcQ/aEBHofgt9km8XvIvP0pqROjwiq7vrVp7ccxbZOhJp
cEfrKHfzxop/HxKbvGg3bT+MVZSo7Op/Z8CWSCPnI9uziMZz2BLEX5VZToWgs981
y0Y9u7YTQP/9b+v4zJSmjowiBKUoAgMzgPe+SlTL9vorLDwsNySc6jLOzjC3S4s6
6DRxqYWuU++ra/bmnpf9e0K7Bi2esF3zJj+tnCEdu54XEXDGfKjXq+D2wZGnYN5c
opXr8HIteo285QFCsGV3s0yKfq14xl6cPJE3se49Ia5Ygp64bYFm/vih79gdsfen
LPyXdgCESAWDdmhgv5Y9kp02oDaYijflkluGwhJBaBkGVSgqIyJVXNEt8FQGZ+BR
5idLjcGSGeb6JPeczIISKLFBGfrwuTEEV8VMotYFD/aHvKYDbpN+yRddCXGO31CO
b6odePkTudRRozoT4+RaDvWF+Aw55c5A5FS+csOrM6RtN9N0y1JnpiHaf/eMeFUC
UENTMnNhca6wPA9YKPha+pVnSVysg18ZP/+k0TaBfUAhVMBfhbWZp53OGGN9CWOc
hjZzAx5oAG8YIVFQRJwkssVH+KDgeUDjkCSo0XQZk5hgtVBqiQeHTIrOM4uV+4U+
sNp321rg+gSi9ZQ3IZ2opqzL6Z/4sOAZxfklTkXi3mpD5jbxKyfhfB6zcU8rrmj8
Tmj8tyFNNfNCdbXEpO9eGql5yqfmv6qxAnJwvvfmEA5UAmDyjQlgh+tn3QbnkPuo
ztCREPzjYXkrJ9OwAaolGLY81L152joqUGwj5VNDq1FNljqVo0Arww6jCHQty3PH
sFtfCcpGoG6h1qdl/6hBY4X8+DEi1BhNTf9gmUvqQB6bS3g+Rvliwaz2hgw2QN+z
OnTDI7qAApejilQE1fG31hmlI7eXuVgx+C9vM2GXFOVfKZyO0QeH+0gau4GTy3FE
NsJfcn54vDhFoA+xeMvezncEdfhE6JUDO/hUO8ppeSX1DZuaYav8Tdp+plrBli+j
T4bmtYDYZLUUsNwSZNKDGGUyjo3734TTYIN0w26XzVrQKok5QECi3dR74xAz9l8/
W5eiJjKwu4KSacAf4WuqaGe++v3hykmV1lr34bsV7lzeOB4nR4f+avXona1v2VVh
VS4VkHxUEA52+VwQoIuIvrr4YKG+JVi1Nf9pz8oTv677RNtzZImN09pY3x0PO5MA
Jz8yiDqgIgm8Go/ALOMpShGSsj4/3HIc0yoeRl2jid45UXtGLrQdbPoPAZNu/Lj+
D6Utiu3gmhE16IKk8qWUM5D2IAj9nAi6HU2h8wulVBLgwKY205oiCZWyQHU/9kzv
f/7nh4oKHlRasNXwIS3XD/ig+YyASRSDqEbkQCYfws9pUFRfq7RrQ40v2Rn/wsCQ
Aji/d3JmTXJvjS2xbZhy2vuBXXDqDA1f6SlclNmW4wmE4rrmZqd82GOylgDMkiot
QTfVQkGuFLfLd/1MvAmKLv8oTAhGTjcV+T/J84pI/NI0ZUXIlFBRm8Ri/T6rAzoZ
bnqIPxMVG0+mn6D4KtvnFMLP3iRafEZrO2Hjnaiu5b2qNM8Qi59KnAWshVpjtMhx
ft0M0g9UZ9yuoE+sIK6trZ3rDmxxuJSNqV0GwYGpUoILeh93i5q5ap2kDUhYNU3Y
2dx/z5x6yLRcR/lpSVi9kLf2sKUJqZZgmGeRwf+28yuIrO1MwES1o4dd029CttA7
BZ+BeNNzEPLw3R8iu/uq/PlC5m+zXwFN+dskPB2G7eEOQQyDFEO0FI4erqJH98HB
+txza7jLfu9i9mmTdUBQOf9Mt3BjnNGMY2Zztd9s4LpuZfkp54q48q/R2Mkf5rT/
bBtgWdG4kG+Y5AZeCY9LQGtn+KR2Nf3NTMg/5aRUkKoX1uK/glZUsvZ+N8zTiYFm
KXJ7+yHOfQl59/UJ5RG7AiHHNWetxRJIss+TrX9vXquhl8vFM3oyuoEMY2X/u+M0
SRSkFJYqoyybfMSja/ttGZ2aaaSGg0en76QPhQnntRWotE/u07OVlHv3gTT+ac4C
Wr5VQ57gZ5we5ry+tF3H7xmZBNG5I74QgBGBqP94OqPpN41wmjzPlonzAvazU+HR
kVjRKpD0HJOALYOvsivvje7S9Mq/mYWBTz9Qu5LyQKEljampVi0ta+b9RU39xj2M
fBSGuquxlkddK0j9AC6qsTPbqyWHK/7ujsz/bepiiqfYpARylNsDFNknwUzFFD7h
l35RUpsi5Z0y+oVDNcXfrKjx8xzAN6VR3QtNZRaDKUOooSXh1l2dyf8Yyn7rRpQ4
y38pHg/DkFAUh79QNqBO/SUstht1vMm7dC8YDR7CIFDoJhOs8Q4E2HlCzinnM0PP
flkpZ58yqiA7H4YDzntb0HtPa74YdTpJnQ69BaUBkLWrE2mlZxFfcpf8UvNguqP5
wRhSZ7QCLrTJ+XeWlRZqWSeN32QJUbudR+xBH5gUXJd1g4QMZqz+/my7UxC4M0SJ
RQMe5VE/kKHIVpdgEZ/2aqWoGZp2fmM4MI/9HQLNueem/ja8/x0/RF+3oxzyYH7M
guMCXNG7z//0QSBBLAvyN9kjZ/IZ35ioSlyx9fS1VtjvchnFABJsE9LHf03xEbvB
DeHqdiQh9uxy8A4rcnxQTgdb50hoHxdPCmdR70gl14pVGwSVimiCMW7AJpho1spW
VF+BfBmhTTg4dyICgxEv3PRLZSLoh1xT9GWiS6QY83ivgA4WzkIIVUBNLUTNepDa
TGC8/ZccPd1nz6eZZsaiWHcQ9Zcp8q6Ur2C2BuKidIabk+fPEJzVKadCHG/vtuGX
WWnaUs5my938+2xS7ZvMLBD6fobPknZbXUn9pN6n2+JI+R/A5TPRsJ/BYnKreOz6
oQ7Erg3J5abOyozfifvMLxoHP/OWpaEEb2elrwz/pz2qpX2dx4oJDO0NBthIkGMx
zzDocaqMXb5+5xBFC62fGGJ1ZqQ99rKxpVaGu33GCjmJgLgpirr/YwXoNY6VVxTr
Ou7aU9cNH9xRQ5k9wMTq9PfUatddm1FefDn5XgntvAgcn7TbIge4eEEA4p/VX0v3
1vrVeHWf+QPZPUkslUfOe8WjU6+INKZuuFkxAYz0PlIXbB0mQJrGZJqA93DUzHlI
SOQcQPhoODrLcnVWMC/2q6CsX4Yw5/uGoWV8hbWgdQ43D49V++AiMUHF1S0xmWpI
lKst8Hv8hU+C1vaA3eA+1RzxNnVSLvmeBggcELSv4O1wItM+VZ9+rQR3gqMqFK3B
3jdLupGTar1brtSGXvemPKPDLhBS0dY8HnZs5qI4TcQ4w2CSeuz92oKCi3a9XnBL
qaQjMzAM1wy8qgeZoFVVshjTnaKKkXAgUcGKwbTj/ei/BzzwQZQf0X7j59I/t/He
YRpWU9rHwv34gOdI3sCUeZmiynk/DfMRtnNjhNKYHgEE1jIt+hSdzmOdAwXmgQS/
WUXN6PYquwE2i8cH2kc8TY+RRZSUMQm23y4d6jb32how+q0x5glNUzGB6gdHl0Q2
UM8rpPFjPmlJZs2BAsvFIjYVjSxjIyA2PQrcMgFl2pZ9cTS2J3pziqM9p9qcsQ0T
8gxL2L0a+9WZXimOx7MUc1HRemajAh40IZnBGksUAFfI0jcFSTzDstM9zO1zk92K
Qqi5eCC3LC2M7OPiRzdKz/DHVOOwuwd8+c6TTl6TvbVLwY53f8u7pLLywxLBDfzI
Y3+u2Rvr9uBKDeTH2vrLhljYiiq4U5VrlnccDlQ37I9Q53tO71UgcxJ4Pknpjnr/
neXtqCo3wDjGOBIyoIiP4BSL0a3shfvAiXnqmR+a0sUXANiTrHPqT8UyR0b5wRvd
ujIRGaUQP09JaP6TWCJ4x8U0O3x8RJAhMz871NbamslcQO55MN9j4AJ2jOqs7t+a
JjRT+r2tdBABBnMkmSFK+xxyXeKRPsTW4AJSqcoL65vOKQXcSnxXbCNCUun0mv3S
Lg4SoJzph77KibsDCZEHFdNpXnI4DYiUF1u6EfieVLFLdDWlgD6F3Sx/m6ipAQme
wxrlUCPyTPsIo8U+blV9nItSBd9L3pfV4cPuoUZOrW0AXbiWfIWtNS/pXT0Pqyjo
QtkDxE2iupf3ASunsXmAle7HBVJgrVogoT5MMDwgplYl0VJqzJS/btK8uy0zmiWO
r2lefeYOVS6e/nUd2psOhZSLelcyjpJYVCTMCoM9VQsFjL4IdfZSYFsStEVLbvDs
w8ixHPNVZL5oB/HDXygqv2/65/3xg00Bd2OpE5amkHqBoqwYL+MNXKsGNf4skwfy
bbUvmHNJWVskByE7cNkOw9m5uAaSp1si5t+5GkwgC4lf9yvIT9sfCUuu7ExHRDy/
eHrw9NZ5jOxIEDTNshmv+aHZJbyR1cA1I04k3tsPfcRmjvQy88com9/H6SUFzcMt
NLMuFLc7T8tTXS5Q4kdFs8joxlFsclGJ03aMXXzEzk98MNPI0S5O6ck4d3uZ/7EY
zzwZ37pt+6WdU1FyhNRkUue0a98V0LzvX6WWSa8FmMgYPOPYWARrEbamMHsnasKI
s9oVZzaHjAW96SfOF4kvJtr/98Qb+p3l9Urd3iDpSrOssCJu0GoGeiFTCq+2q9NE
El+bHZEUSGYxOQz7e44OA8PQnet/YS5QnOTO2DEhruLxoEn7R18scHm+SdjAc2+0
xf3LyzIDK3AMzxcBCDkkwB6rxhoz0TOvW1OfOfCHuF2wPiAdi9NCfNCUZzax4ZCJ
vguoRWesyAY4a45GsQtKRjibyV2Y+r4xLzb+oKioIZXjRvJNGyrL1HAL+QRDmFxf
sUHmZBTcCdv4DjNdpgxC7erYJcOUJT7mJPmYBBAL9D+GdITEb1oP4unNpaUC8hS2
tdd3rkCHsnQQH88bb4gW5F3Yblt4brV38s7ZT4RM/sYheg9RaCpVJ+4U3GfhVlkj
Vwi5AXPd1mZzoN7Hk/DOlPm+FYVYgRXdJf6u8q+4rKjS03L7HZE+ctCoEuIbproB
DZPzx8nuM57h+shuIsdCf1+IPyCb1kzXkM5UxjYmqJBSxfMTB7BP9PlV5LT2Cmri
ajZw5uU/LviAlQmuA2SX4m4woUOmtfsfVK3rEDAv+7WZMZqkjvYa7MSwiZQvPYwI
lyOzQ5vIppML48rSdenNZhjNQvdLRuGQarOL0bKtVblkkPh2GJoToMIPVazhNXKk
bk9Ax0WmsiaMTjw0puJTNHZQMbUEXV1/Np6f2aTytz6KqDRctawdLUCC9F4y1MBX
4tgNpRf9i6R0XYi33P1rH5ro7zuW+N02AfbsQ0LUSYaywJ+9FwWFWnuReTo5y29i
7VMQkZxq5ugw9Xpky4IXMFq6e6akyMmyK7tQGZXRk1ICPAVTc4rDWoWvF7TzV2Z0
QnUvvlJ1mlXCi0VYfYDdowEKEut+sqWRWjYVODPz35B+21cfd/w0XM9eGLzEDprV
bZ//OVsxunPNFUN7XJeomlNQJRveTsxsAjEghBvYppmkkT/gN2L4OXl3FodoQovU
1n9A4oWzjAlcQKgvV8Ht6ZqNWNFRreupvjVcWuUzc1ejZ5pYZi3wCbK3zEANnJjR
A4ObTON5cIZOmfeoPiKHxJQ4yFw6Ob/PGXAY/Eh4PGctmzh5yR9eHlw46iOe9EQX
tgdQsQvUzbz3z6eD76b3/RET+7L0RRppRJrbfhYekRJFkK7i7XbonwAeLRKl3wt7
twtd2F+Ya1eVnqTsmr0+uZ3us1t30/V4t7jPPW6TUzl8SJbhZXeQ/PPyfi4md6yn
fXMOWme1lHkJ5nrNLrHtHpXB/2EgXGCbHzU1is5OYNA23GtmJnxzwSy/zmofFpUJ
GUNDe9Nlp1ApoeIJe0v35jJr8V0pZS3hV5FpICzvcnspKe9MODzQF1AgKP9UWVpv
bgXh9c4/edgsBsAou7s/wtwfMDPhSzV/o4f4x36Iv+JKAPnPvKPmbetYc318zYqW
LLQHY+TQsW2ZzZIlmYVSBqpf+5PexsNfodemJMibBMr1OzhWaPzN5eNfPU1rn/P6
8PROPDl4nrJNoOAoMXLvcB1ClmYz+fGHFAebR7ezUZncHcAfhcjKPDHd8UT6THpL
uiJuUJOn9xb0uKaB2p/AwJuVElswNHM3bq2ICIeFHy56UlIEhplQqnzeDThxC8MK
AnpQK5BGqRiVfLRq+s6wzYXdx9Mb3+X7m7FucIJfzIv/PYxgHNak99HPtEobi18E
9x+T/3PUXzvDKyLznbY+/tOeYCnQ2mtVtt+v7eKOB2cc3SW01QzHqa3YpLl82wby
j4lvChAnseUjvG4mlLGCdPdUXuoha62FvVOD+7xIHlv7cQAP0GbcDLJPDzncNL4I
TgO1VXQAwaabvQDzU3Aoay1FtTbseUDZLw8NUgG8un3SbQfNGQkbIt1ooolhri0B
UOEhDRO78JLps9g5+YDO1HmrWSbIK5WVkufPTV5sD8w5UxHEzTkCYa4yUVW9iwwE
3lBwpcf1PTz3FIkbxi7/zZ0d/NGk3SWAC130pQQAV254qT9HpEdYUyktkezCWpXF
CQ6KJO22B+TiPas810hRcEuP1b9RkBocrjVlDLN3rBSsejk4gGy4cjaBNN1nQn4Q
L4u+pFw1eXShZX4vegjTvwMQIdESVrXIyONg8S40kdV0R7Sn9n5abTvDHjTjTgV+
7nuTFAlf5wk1ykJ3HXCqpwXEK/DeJ6QlEwmVtIUiB562PbiT/OIiSjgr4t++brJg
gwylRCFnyLJaBX29xyMlwgCYV6F+hlwV3hyNNJBQFszfL75YXmqFBR7kOpcUDuG1
73Bco47pIZCnZpV4+lwPJjZHZSH3n0sCujZ5fHPlxdGePLA8jp5jWH9NMGGTmZDg
sM10+Xtwfh6oWN+WHbSus4EmxE6+yEBdfhxaHorPYA7AMDBr8v9mlw61jlaCkmrP
++NsND9xhKSYmnVUGl6SKaaQdZxcflNYp1Y3WkeUoE5O0UNsx8GeMLcPQqIUvill
6SwiiC9FRtw4HgWvH2eQGW5qXKpfSHvoAhcIcBsp7jCezk3/3lALk9xRV+HmU8R0
lpcu/kaki32xiNGl9+9cJMSjNpn/Q4b2QFgkq9rLRxpQ4C9cU+Tn0+LlM0VTctX2
IpW0JobUWLM7ZYWhVYghqFSZMaI8WP1riyR706MovzMIWAmsi2fiLTwciB6PfGLh
PfS0nh1vpa55f7p2uxxToNKrUUoGRIlYApv2dBNzgWC/qJOjGcA5Dsu28wbD2Tca
Dq3WletUSmiTxR3kttx5p0QmWqAdbCVIc3dIXgR9OYphaZjc6DeBwFYJb7vi9hxW
0BEvEWIz+7l5ki3OZ3SIB8RqXbb8xcUGj4jtmuldJqZyILtVO/NnLko8Q/wB8/Wn
6JJewO2/FXZECROuuxS+H0Dia/DhQpANlbziIQ9B0JP/AzXdJuL6qeFHwUNFaM6m
MB/y1RLXiGJQiYcVJYaP8hLur1RPcM9cSqcjGfAXqx4i0Q+zyukUFtbqkgPAKJoy
ln0feSdyDEDHO2zfFCLyPH7ughZcwQYYx/inRPk7mJH/eeBP/saHJ8+N4UafSvwz
4Szwr07z9rQhbR691Qkj420/MKN65qvehA/9UT4pW/osW7QPDlgVHxTCgshjiA7+
jmDDVVBsyIuFhVoQjgkN+M4k9mHl/xRqQsiWyf7faWWZHgKx5OZAbSWDhOhL6OPK
qp3T/+0WZxvHog5pZOWL1Ww5Hxuf9gcWdrUELzMt/4IE3sAUD1dFmAwjifII5lVi
YQVS6ycWE+IYT0k54z22yJlZqvK+AAAOCyidoBWNM5wATYvSkYtzEjKtFD5LKkxD
yuHprM5096LgfXLe8ygFWt2vt1ALHjB4JhhsOXR4nyQwzfnfccMtptV2LybK5PjL
tWakQ5MHBRMXF8ZFJSkYZPhPIkjlPyBXfXNihjL4Rx2PGp5+yNLL7jIkpSQ9C1pP
HUhC733xarTtzKCtRO/G2SeNG3p4OtwWDtxEfHj7gNCKS8QG9xgyKds1ID3mu6CE
moVjgHJ/xRAECxUR/+xuXfF4CGOFnJtdr8PJUMC1z3PyKX4/DqnfAhyizRNfMJpa
S10OGVoT8kcD3XtlrFpvlEO1J4iQwVrmA1kXJ6lZzwulec3RG/lH3QIpWZUO5305
2teSWdlDzgoD2/Uwv4CnFez3Su6oEqWPTbiS78m9oHW9AuGQzUxn4eA3UH2/FjwL
qPpz28X+EH+LSs2OhArbewOTzD6OXiuG7RO1OtHnEhnD01IrEYH1VvaoNmZo3/dK
b82gwTuY3IRb1HS9IEvdXz8BFNZJJM+s0nsg8m2H2OCjNFkltMm+0F5M+DHsFdSR
RhCALyxwMdOUY/Dqg+pQZNBYh7+ISLdhf194JbOF4nzt3HGrba5d2O+BZKFWgjWA
/y+spQzFfGt0k2Lz84D81Ej0O1KsXeG+q1DSKZhpKRfjhyq7DpM9oFMqN54myIKC
N2OfZwKEivaVp0juP+APXUhTxizq883FkQsqWcQ90s+afBPit6QW5g6L+pRxnTrS
QpT+gohab1blkDIKk0dTDOwdF75OEDn2hK30hGDcupGCPSBtjC+1/Amj6Zx19zIc
lmtBHOZxGSYtP5bRCv0U2RE0jYQex82Bsg+OkU/oJvHI5TXmRvQZcFmhmKzkjgIi
CEApuHptTua9m5qJiPHt5XDwLBns9l9X7i/yGw5+SCcuUQFP/pfMIPohyk10W5Ir
O77OMUiFeJ79rmFBxSohEF8FMdDooX62WxBHIIPiMH9NTzFTw9qG8j+svp9gYknD
4nhUx3pwBsegGODZ3kVQtlmQp3Iml+G+sW/NyxOnIfpL03wtYPmoogVew8ZIlJ9O
oyAXqpbRGTt/RGmH84lcT0SNVsbma0JKrMhu5R+gMTz0GnEj2LUin6l3BC4etcok
xzsukNBnvel9RvPj5aSxlL7zriQet9EVK8b1pEK2eLNIBKcVqJhQlRzMMUdPwNUR
JjaBsKAeo76JpBTXEC3maXqFk0PH0mAtjCJqpwxdgIEC8oMEDbSeCr6YT3WNNwPu
QHLakH2YLo8ZRG2AgzB1Jm4tJ+luBo3LWqB5m2qzPOKRGYP0QsVUAkncCr4VZZy3
4wuhvGJxk9LSYZJgMTSSecyiK0+WanSPIYTWmsIG6nc4jjX8QgwZ/16mdJhC47nw
MWQMp7PKC3pMCzpSDY5SuAuflWNpCSw6MBF4q4TUIH+FUZ1Lt2/un91q8XI815Dr
pVyks2F2EXwwULFdVSKZg+IiCRkv1BzHl5eq6v3MIckui889FrRY9dw+LPLgGL4c
UDYldoFbbe64xuATiDLp5XG+7KqhdnKDGMq3znTtS8iN6FzbcD4+sRmL6bRP3I3a
0yRl9JPUieZJ5zd05x2GJuYWn7PSjsf8E0B4Hr2vunwwEOVQkjPsARCXnkrRmcMe
Ye8wjlBzjr9ZuZG8+/qRMClQC3BDICiT3SIUjQQODSaTbgAlAVBE1RZclqHPL+ks
Qu4VxCLM+XXnWI9HxdMcyDBqBqEu8rOLsVADoz+96LRWOYcEkJ/4OgesdZxMr7a4
CY+rTASRXX1K6U1tFAx58+QNoxMWRZAG67IezDoQgh+nQt1wwUnweOi5ZtV4RlUm
ydvSSvRj7EPGuyDKVJzjlDQC+5tE6msicpLe3fwfxqHQFAdbgRk6Kl7oKQsHxws2
Vhdna9j1CbE9Lo0JBHW9088+H/dsuxdcCFgwcSW5eiR97YWzGVWOfD7f4qqF6rjd
zsCVTsbawgWaemgM4MgLaz+N7Wu66CbXnGJ2fHJ7cBGijN4hG8jFx8KTySJ0j4rl
FGdZlDA2aPO7p+/roknT7XPeSa18+c2WVjLVOVvU7Wczy80zS0flt0rgjSHkMVDX
sYYRZPnd/3sEfR/5P7lGkShfzDBWaolf3ESKVTvAW3PgHZQypRZCW4tISmMmNnmq
2Hc61EB/UpppsvlpqgaIC74w3wj+E0e9oeeRBVCMINtof0g2kabyCP0LwYxMGX58
olQcig660DIvQEdzDDsNjdm6HGw33eHQqyC6TuHBKWYZgIGtS+wdH426EJM9I+J4
SQelrYs/f7uwhK7XVdoyUB+XbGTNTc5C8tO064qiuwPmiZJkYy6OFlhdlGmpVqFQ
TwHOuVhmTgIFKwj+EDd0Tmq/hPx49dnB0Ho+VmSJZhsd+RnggrLmKD2GPD4QyRGs
fHP1pHblJD2iagCwaEdeTVoPXYZaJ3XB+ZCZUhjgExBhs/iuZjLm85NuoVqHjFL/
cYl8aolgRQe7pPUG6WLXTDvi3SHp1LN+dnrkFA0/VDSQCpULNuC3nHwEHG0MqLv7
fBjY7glH1IxGJ2/KPj6gOTizrXU13kp+I21G16xGHz3dN794d8WJKSBLPIYNWR3+
s99r8Y6uv8ow9A+rZsIPESE9s2RFgeQReV1E1hvXb7niLDAbIeFhDuKu739a/ajH
jibJzxtjV5nIC0+y7Z7WvpAuSZnRkDC+jKwLsjVp41wTCo8t50f3M7K0yZwGghFS
3fAs5at7cHeB859Kpptx1S9KrL2q9jtYRX8OtnQ1IwvizrsLAeU29/Wu/wumHLgc
0OQHRv61Vh+N1n/Sj2feSTHWEvRsYrdK5DtWQFxKTiaKZvg3e7eSDuYpEqlFBU7U
6eMU2wyNYoCj6xqPSwCuyoB+ZF08CgWD+ac/yFsEoFYAonPur21Ae6JYGJLDE0E8
WDQz96l5wKppEB4VOzEsyrhAQ2sdrGy2MT1wDOTpLYP2Yi6s+3aQ1KaK1ndNPymU
KHix4fSnwC+Lu94cbM5cuTpBKB9+loQvBuYI1kNknFPYkkNU2etjIFS26VWC6eAG
8UfZXyHkN9pK4y8onn1XivI+6Jio+Zd9L8QPOeItOVHi1NkWYMsLDfOOsULSkaaZ
FNs2ztSgqZrD/OSGF5JVknFswlhBzs8mfvxyWGg4npj3hibUEINkJVyvK3fq5Gys
H/pz1+wIqxtWMnTjoIc6pfaCVb6WJAUZYRfbPbR7Tlg+2yjt944vAXjf6XioknDU
bCKJKwoRmB/5S5XC59xzmwKqxzrgVYlCHPokbBTgnmW8RMTTiw3yCLMORcaPqCcz
qbOLe0YvYlMGt5CaJdx+oDHoqGeOxzse3ogK0WBMFeEE2irqERsf1LvIXM0p8q2u
Ho6mt8szThCQuB3vAasYrUgmc3gPLfM9XMUrmDLc+r7EVSt2SNFrLGwREGOTVfPU
Aw+H2D6tl0d+svinH8keBeZFG1ZRFfP5pX5V940odc+XhUGW7UMQcKWQobrpNSoe
dbX0vRdlae55qXgOMaTWjArKu89bZBRg/+kXPFKlXRzRVVGAiG6tICR8bajIe/Nv
N7sVXrgbZoYyRWQ7vFm9GK4bpVlWqE3YX0u0mtJ6jl1jJQrf9Mi93ne7+g5/9prR
+wICw0gWVNjaq8NnDqX3wr5bga1ih3Sg4RtnUVNbreyWIUrOZ3B499QNIx3hSaDT
YA0dXpp6fQaZpOhJSia+J7ZMrVtyKvBnbIz4JoKfaDrvyvljpUQ5mdk+IrJx5S5E
3WUzwEmCYkoItDKMOWYhfnrwyG+9r5YVl97nr2Aui8Gp2kNOMWMNZBgm/fvs8UEL
9GvnUwAbsIMaP5z+1+X6H7sttIWqyM5L0lsOHz3Q/Y/mg9n36H0X5wPznY5JpKN7
Psh2beq4XYPO9b0ex2hlYosVlWCmSxSMIfcRu5073TJ4I+/NDfij1Wt8WdEAsS+B
OiFJMuzz+cJ3DaTNfflmme2WSPfO479UHWojVuyMGoQ3aeJZ+xf/JCi37w02oB/+
LHegDvbIFMUW86dMQda4/ErbmEB6DGT0i46dKJR9L13eS3NnEb6vbRfqbAlANTfh
mdZchTukqXgVMdijwtRIgKNmDdkwoGuCTZWOocdKpx2DGw1RNRffRtOWRTtWi3WN
3rbKbE92E58eVFqURAdc2opeIP0CQhEnLfaCx8sYoKeCfN8S2Vu3kdqOjZeUoYg4
9B3ieOs49XZFuvpu8NbVhd7aFmdwduoKpGbDMxlFSzSCPtmLmJoKyxFeFOsfbXOs
I+z/pxa1v7NP58AM5qeMhXOv0+MhZQY4E0UStCbALlvMdGab31n75cX7yX40UNn/
Z3hBy3gt+30RN0ZdpZF4Sy1jkLATKpLq/J0aTpr85W2zjn+Z5Q3V51AFQXb/i2Hg
3+Q5OEXkzk2ruF8NG5otYB/50FQ57Z1QSeecWANONoZVSYSodZRC7gDWufMJs1xC
zW0dy82K5AmzXFrmWfWa23UNubWlZVi9CN0GsDvdgLvAU2YcD6F8c1PpwsMgMAQW
lCXIjBv0mnUku1eKNLodQb7OSki06ORv2NRWngA2UzJKO0nX+J0J+bI2LA4lwW74
AMYxC5614vhpTnFiHl07LjQRHDf4I3XmVwCTkScq2f9jED0A6U9hC2E2lH+0qhxp
IlrFkMoq+kQ1v2DYiFyM+fncPLD3QY8AmLKiQAaYzhxwAtbrubegFfRDgesIlWO2
3fVyfUoE8vzDbzDm/z7lKZ22205jIuAp+3qSBbP6KSGYXKt0lSGUYCC5wC5ZGNVn
cq+PScZnhNGEh7MgNCR74RaPQB7YY2LFhASxRuRpTRBA96stmLAavHXAeJQ2QqWh
CpVBMpl8M6CaI5ULuDCB1Bqb+ux+w6/78sTvBj2yA60yVDCc+kkq8bbMWbQVmpLX
rwah7iZfTHIYZ3halMjGtWqqfSTTWNGmMFEaVB75TZrGA8iEi3plFTLLO/qNTZlB
TkYJB4CKZ8YJu64YPqtoue730CIecIvsjcxPEUcCce7SuEHFp8yYsv/al3JhK0rp
xzG+YmLMRxjb2nrB3oaJ8fOGHOabnhMJEVjUSUU/ma+s5oVaBfyVwsafjCVYp6f8
Hwln3/sabvAbBThV9QsNTTNnRbKDeWQm6sZjwtEJeI3ALxohO68j8+rA3x0dUqzZ
7nGdBwG832Xe8EOkDVhh21bcNuBcEm4DEE8iTg1sy1viebWCi4CQj2A1BZn4XAUR
iuLyeoQHF2mHMl3awB7XmrBMao1auIELQWGBQPllxA03XlEsv0bWLkzcFrZDikYz
3OA1+ojaUerLCFwDcRl6qzoejQojXAcvs+1NHonHnta1BWnHpp8BmRABo0d90n7P
mes7l6Kx1bPbr4AA1BLt21KEzoypXRmTPokjQN08OdIt5b7/UgrdrrKjvgpr/SN2
gmVVpb5vM8kfnfO482zusQqFpr3xe18GnMpOluDwO/KTsLnaiZRC1iDJwDbM50rD
8wkQfGRDbCuMJctdkxHAQGlIRIa7XFEAL1bCzWQ2K9dgSf5ysqkuakK35H2zfrXV
SunXgA5vPCWqAprqg336g9xPY00cy2qwc6E0Rsruz8EDmIN4s/lbgkkxjpeoWmT5
I9VR/SD9Zg3p1x5OkLCXZRDuvb63VzxHLXCV630SnM3FLoI1UpY8s13Ff4xjiBm/
MDS9gJVVLCp5CZLQlTklktAecaKSjVCIrNBuiTdPAFJH+IKEyxViHwAT+vlBg6v+
AO4K6+yszAK+xgw3Q1Xl++y46549NkhPoXonny1ObOkUTWBSRrmixqKvSLndV9is
EyuERiPXFsdGUWn8v1kA7Slh0JbqLhoNh6A/jXlQ/DsUS0KRD0t0ozuA6t272uln
lIJvaVu+XraeBCWIs8pMnWX0a64HFsYZdPzr/WV6y7w8jbggOo5X8y4UiZTjF4Xv
TFaRZfqyPmqMFK3zbAGzwtsB0g+N8i32E/vSv6BPkSKhwsWQBRt1VNwNZMG2sUNU
PF/7XlJMYOZhVuqAIIe9+v/MX2rHvDRcxezR5dtI10QBe0WLv74fTHaHyPGMTqyz
SXHoodWxmhvvIeFPu25VZVe3s02OqjwFOkVQj0N+T+v7R4/LOe7xbDGCWGbm85bJ
UZEvbyWywvmPao/YhhE/ePs/w8SigexPXZMu7aWhmdOmO44AfOuoPvaVMFca49Mm
rgiKUWtafgLXNTRzgpabQpk4rZT84gqCl6swPEKCQCCaHx8BvWxiFcQgGhALACd3
yK2MK0crQaDBoe3fPXQC6LExw9qd4vGEy+UKjH6DNVh2bVopNBe4wh5IZaJ8Ykxk
hjrr47chSDiyiEgE+RUuXHSqDTdbr0E9RP2jcjJH2JsXBptCOurL14hccf1Euw57
WHBnYwUAsyVIzcBYXPqLWM6RNGIrLkxSAUILb7o6pCX+8L/IQH0ySvzbCJKxeI6h
JOpzfPSJcdISXLW94Ydv0s/mPYG50nNxury9wJuFH3+5e/PTu3i4JZPMQJzemox6
4rQp+rdrz9PlBl5r5a2ZHw+mbtLBfgVpjnpvbPdruIZaF/SKItDicsT6LxOlxkvp
jbpB5c37O7qDauPrhVifRT3a4Fe+8F52YWHxEcuQuIEptiyk/TLmLeRH1wVvUF6z
oaQIWyd+nXs8FvTCcCXpA3UIiOhAht5sC5z3imqp2i7Bmo0XPSG/Wv0aBvcQ2upS
Zesp0Z2kog5h8gBR3s1Dq0NZhmoLkf+vbVh+lIzSKAhj4r4vIdzxdwsPPuTmRU6V
wNDKN7wlx7ceMSNNg8jRpqaVnfHCDrsjSMvsmi23WRhCgj1PpWYtDUcE74IdTLRH
8IJH+aLOTLJdLCZmi4l+MofIBkGILhzgLisXnTkxCFb8ZABR15WxSrJ8UZPJuGdk
QUJCptfBXDiASmcc1buEjoGqSR1vNsogqs0AD4AeCdovQAUK2wxYP+GR/ymBQmeZ
d9pSjMePi45J0VJT1XqfjxQa0OOFfpsZx7kiqCGPejoa8gnOcaxOO2TKNjBdCHx0
08FSJnUgIiCh1+rX+x/BPWi1d5ZiwBSdh8k/Z/m8vENda1aCg4Y9SFy/NUlVNJFH
LR4j1EhWVPf+4LFLvYCNk5fakOF4/B/4tuWn9ZcLt4G+J+bpUOVv6G3zvUNCl+Jy
WLzjHHlLs8rdy15VY7zJj8O3/OYhcn8X402skkLpdGiHVDxyMMK+foFH5mK8w936
M0t9+j6YFTmySOWtpjqDrAVBa9BcTg4yxiZ3/L9UMtuI7BBUBU/jLHQoN1SSIrgl
I74oBtEe38aPgusTFUruoz+6mK7O40Fw7Wp00jTrZe3usujteL5GsoBGbmpuU0S1
v/bRZ6Z14AcrzdedsYuAzkGZa0y/GW8JWdef3T8dqCYfBXrwaANZoThG0L0B2WgQ
GaalbBimJIIOJ+ya8edcnUxpMyJiKlc4cPzRPP0H1sXkk2e+ZGzzNPAvJz1O1QWT
Wo7Vzm0NseVppqet4bFpfZrFfAps1KPB82VUkcIQO8cDJUybMCMklGSSuSCBhGoO
CcLwgo3QsQGS0X+qSjmHFwhz1jAO9eiQ5X60oFmgWi5afNVXfBgj2wEDVrXx0mAd
UutBdrMAjiDo4H47r/VefGvE3iz1ZZ0VJWb7t33NsyddanofQ7UZHJ3Bcr1hlhPt
Ffzcp2/nmZ6xgFXZPrSz04o7cFacfbnCE3I4ToXp7Y2ynsNprmmQ+jUfDbA5Tqhd
dU+PT1Lpjxum2ILhXm230Two3FApgzHBOJwrwcCsSuV7qsDwSmG83iilyVHOxOcF
VY7QfHsCcNvrPRVYGaNb/Oe9nrK6yiCLsJjq1SslJcncu96C+2tKrr8VhOkSt1pe
OQwLW6AK01GUPnUyyu/dLTexIqT/2K+MrhOz/GR4PXBlS105iS0DOB2LB+DVePOF
ZS9rMffo7hB0JCtCTQ/c0WAJgvXp+6Y8c41kHJvKV/2uaM8trCNkBqQ6iZ5/I+ok
fkK9EvC/HShsYXZont2F1KjYMp+/GkhEFp48pfaSAqYXDa1G4bfN49pffsrm/Rtg
/dYI6zxUi1XDRdimex7/1cQNqNxaJcd1tLbGVibwoxLDQNgPFLD9HTmxrhjiGs7c
J4aELrsFMG7oFgiwkNnOsn4vhe4E++CBNKx3zTk4UQR7RisqErK8DIhlnvFJ+uBX
PzW7/Bgm894sOiKVB/fKwZmzdKrz1T0k5n/YPYPAbHy9vHzINLQq+bcvY4HZqyQ6
n19w792pRp2fWPw/vmy1/CorOcfeX7JM0wAAlvp7rgTdts9mrDvdgA2e+oCbY42m
D/J/Y93KRI85ue1dfqVqP+Pwnu7VAsl9WfZNPk0XQawq8RKpLNy8KKoWd4yVHjDL
ZWBODCG6IiVcMoDzEg7/8ND9NRA3PS/PrHt96idPXB4V/quUcfIPd9h7zOm2k21f
TGoYZOaKXowfjZEIrdHKjmI2QNIqqJCUjqa7jE6SW8AVz/Wgq87M7PTDtqoQMp0e
KHteFVVPXuN3FXmZntYoGi1rkK9/9gYp5wnyK9f979GO+7QbgXJ64LccLPPzwyN8
nGIMb0M0aj6m4APILdihz4RezaAI5RryrFh5KytmXfxjKQl6S6Cb2IabVvCG+pty
TnKXV9lMkjS5DOcBG/nOT9IDa5CMTTq83Uu4jYAEl2TEY5kq7HwIlpa/t0t4rwPG
/c2kvQYWi6VcXroGKThqUh0LfiHiv3g4Zhg/L0VeJYmldF0PhiCpUGyW3n6IgRnl
i8Kffw492k2gFpNkTso+DdJs83S+8p9b36aAPK6Sw5MKWyVqab0FfqquUU0uhQNx
sc1DG9wKef0yJ+CaQCvtUOPPDuD2OwLAOybGHbVf4iahpr7VT3uxJHLIKH7aNaP1
gkvy4Uc6b7GOKc1m612Ojasw7Vu8sXdgg42It0e+l9B8A3pByT1ndbmqDjVOcUGt
EScIZDRFORe2wAt5Zn4VuLJjMFyKiO8JxaVzmXizUrTUbWOTLnzr9YvYR4pvBWzy
aXVgNe1Sf8CFMVimojgey0iKXex6WIAEXdBdldSFtWnRSCW+U0hIaIJFySO5YNYi
yen8P8dZ2OuXq60V/5oPwHax3RczsmsRVWRGnBJvkAzQ+e5VAqf4DmYKiVXNqWpb
6f5qy0U0mfxmkZZHJgKi+7augn3BswUhQgdNjnMk4YCdeqmktY2TuUhlm+2fEe61
4iQbTUbCA7tz74e2AzIBuveQl9Q1zH9n7QrD1QGq6HmcGl02m5IUNxVX4m5kzHY+
K3mXY5pvXBE9HBO0hdjVAsA7i9EUi37HVk4qPNHSR7BmaU9vMgrCBoBquDXk6KQd
Q4t+n6woFaiuEa2t0v+VE09kgXWa3RAwocfi2f78px3AuMLKk44L9QuSx/GvGgOG
xLp3JIyWXAu4UhuhnSQz1rjNJCzQgnyOooiH9JAESvB3UHMMRvfZ//q5UuZWT4ms
3nbLrawm6cgef4wPsShBYEqYSObQtQmZZ0mv4KWA9xFpGvs5Ifmrgs7/ADqcn3tA
fBRaHHa4T/9w6k69jGZRbWGCpVxbCzyf7r++4RRUB1d8i7IZe1P24G+GQKRSC7ac
g0PgPeuIZuAe5GAyLEs+FcPYWleaE/DOrkFrDBMR5rkYXf2TG4l/kczWUkCk03eb
jiNH6UPFKHvREGvem98FvS2Hc3KHzEa5e7pegReIR2Icfne3kZLOFK1q+/JjubnH
hdX9lrHJhrMgXFMfNGLi6R0CzKEg+/zk8KDZRwy4aqJAS7zZJZ3XYdCnDNyvbzeP
VcaS/DFraVKyxXfTRu+Qy1wV7DPAFHpFl+LiMVI/2Yi8F85Y6fYiVFxfKeldqlxp
ulQndwtJ2iglOdsw9tGhHQEJqjbdQwwoafKZgGRRhFeinbTnFB4dAzoQJYfRtWMj
bn0VxvvGmLERF2DhA9My5NkDiDOBI5z5PAs3Ev2PhYBHvYfvnRrBJjRzPtZebZRU
bK1hqws0WJhpFnTllrmEdwYkGNg6X6bNzb7ggUNkEYQcomNz7OZx6xA46eUAzaDk
ZIN+O/mpuv2WWIxbuVVUrZY+GZy5jJ+UiIijNtLjh3rRKoBswTjkXGZcvLBDXIVc
2DFpMtL/mQN9ALJV6oZNR6PUS/zz4GpdO/mDPsDw5hmgu+iealV+WhaN2Ocu5gQV
lXTrct3Qd2F1HS16cOS+Wz0S4+CgdtJkbJXs+r9TVxKtw2bOaTKK3RVlfBoqyoHQ
22zCTjWVTdCmwveahkOJsUhGu9yNqbY+D6tDbuooL23Rds4THGz8lax/WGqh0mcM
TY8DTQQnC58yPBtmr3aAfdge1Sx7EK/Dw0RWfNoSMHaJ7FcABnnZzXRPQbeRo1HO
TjsieGDzjmOBguiA2Bz4jMvY+7qews4Dt9Xu2nO0m+fTeGaEzcYzJGiuD7ucPECL
yX5fKjJOAsn1U1PdplQ6eAa/mxv+NIErnzRqX5Cp01WF+dvXTxZjYkmoH/9Szxr/
PYBqezdII9wuGuqRPcMG6c81a6KOUPl1at6LxGgMsaI0RaAYMDhStoYFsA9IHEjP
WWykTH9P4OhdyLh+QONA89gOHNzPNsqb3WbIhDk3Qy/AzCMiOTEvBmMU13HLSGLF
WsW09q2vuNE0yDwG+xOXAAURqpr6AHA0jLiYxie+EpUAWVAf3hc/Y6zzx88CFuAa
6AAT7y8MMW72lgo+U4sG40cU5KSNUmgP0pJOAUoVlAyzDE0h2UKvaVx7qSO2yRxd
gsJrA9SdLmA6XVSy1mVEjMyw9BDkfNZ3nTGAyBmsV6mqF6NwctQ3IcDuBgwiozfJ
A+swtsYnD1fn042WuszTGeslg7rXf613Fqwzg1RYc1R+kdy7tfl/PggiVZteJzFW
6OTa5/RKYjuy8S1zC5w9e54gYLpSP0g2U8dhu5CcJCqLzshg0v3acz47rggNj4V1
LQdIWUpaX53RTaUMKjXEx7yzeXvibaSD0pXgDmBzc47kIJvAv5jVKGIOM4smRthl
RFfP9/nqzlzRsqlZvVikNAKhmAiDbJAbZVt2ODER+TioPLXaS3YVaIe5TIep8wEC
cbEV8dZykeYcRmnZQvXBzaqfWRo1OUiHazXMpaFLxZGG9broqgIh2k/EN03vXjyy
IN/GekuIt5Ghl7iVUvsHJz7qNPZuEcemR9ye/pkMP2bp3BAYdQmF8LoFTkpdpyO1
Df95z4ziUYwA0qfyNZ0X2BUxfs+yRz3T3Oa46ewWQvSxp6UdTbQpKzowUiyQImgE
ueeIFZ/l5tHE+IaUgA6rqQF53wUmiMo1Ouinfs3+pxS9s3e0oTppKxc0eCHHKFxE
VJ5NR2Z91x7ZBI2qr6KpnOD08urSsnwtYFq6DXZpDLRb8S91tvTjmXGsl/jiGR56
bA+/t4Y1e04L5OSMQVtioktYkNL9V2Xx3H1vQ0Vg/XUPU9GJ3h2IzIz3x5eWpkeH
5unFeRPy/8FYbztRrpQmXMiuW0vqi5DYLIJD+xoGTLMd8U6DRQujwLin0fQvb4nr
4WQdklIPanfKRA7YtGAlOuA7mMpelL+FbfippE8d2PPSo0OFVJW9jIYnJbhJTkmG
FjLXwJKgN4O8WuQZVpC6IuoQdnnQEcB9nqsvYR55c9kYOEGWo58sQIMnY6NdnDGs
2eiozY0emP6I0yuvhhP6PtL9xGOI9UeuMeIoblueAu14lQAkCDJHXwy69XNuGyhI
nSCHvjL22PeS+f8r/Et8ooUphr6M0FXqoXk46iYsUXsVZqts8N41GiBYzXmhM20N
d2f9D2V0NZOgOYMSyaUv8vEcDEt72iCLMZJgzbiLYw9D33eGsxU8w9RjWudSNzh0
i1A1DtokAh2L2Dutd5fFogeE2NWZj/sXXKlnB4b+4TrGfogTnhJ/sOXDI4ax7oOc
UTuDBQZD501u5s6PqElbrXvON1xnFTFdIpTqjT/mtS6O7x5oDcPfEr6WGEV9fusL
59ypVrEZkRIRL1kt4jF2vn2P0VM2b3RIje0rQPo3sH5YWumne4XGryJd/URZnFNo
KRrwcb5qUqRRf3Zbk4FEurT/861dz+tQsQx9OF+1GqDL7cVShJn7WfTiNjuVFHHO
rllJ25tgd7g/7goJT4LtupGiY3l8cUrSVyndxDRG3Ak1tNWHXPfkMM9V2nCgB+Z2
wER33oP9ixjUPzdr+LLC6RkTJGlFLeJUKUdIin4ZuL98oBR2LWMYimOsgDn8kL8N
pD2i0i/CV5O5wUqUwRADGoPs1t+DIczSMuY8sJQ+riBlVn36Mx/lFXMrWGkLtVEz
rAzWps3EYJmO6RZmp43FhX25GoHESSsyLyzcwR2ivC3JxQCiborqESZ9jCi/zI49
YrUKEiTKoe5kMcifFmDfzmpSSKd1hJwwWPl4N2uw3A/Lkmc0OHkFvDgdxoTJaa3q
Up8rAA4uBbl9tALKb9puya6Y2jDiWti+b7+/TCNocMWftLYAW3O2LlEQfvGmTfWx
9+vKBExR5h7+G85LGrdfTrlRNztWVWg0J9ZpCDLM++wui+IawbrCtAKIaPYccVu6
FLvMwzqjCxn+q7HMGFOuk6TAU4AnDOFwCztZnLbKVM2DxgIFy/jVKaD3y0gAYZ2H
jh/3wmvG0yiF6mYSN4Gfo9EV9/Up2YhLOKSIJ8g1tUxaKNZto4c2dRg4nD54G3TZ
VwXvI9iSNeQ5tj2R1MwSg+FlSlyTPh68VpUUBxM+o3QU1KTK9OdSGh0RRqxkImUL
hL4o13EJyBHMpkat+mm7yAPg7uhEBSIleTjsyHFpQykYOfGU2WxhttBJUOrjpLXd
1qfG3Pk6pKy7oP2TlaiYmOgwkIkNjsjedyvAk2BbSfm8EFNiKy3H2XSywYZhYhcp
K45V5MkRF5XCWEB4hotdpOTV7wYgZQ2nowKfH/v8T+jRdeMlMF+fFAj06Frp2H2V
kfB3JUphx1EvGNE3B5F+EaXdoRrS+8A92s9Sx8O0nax52Zdh7TUQMS01DdOjwqpe
Bz0PZwo9Z/dC6BY5rC4pcZaOZei93AAlou5H6dAdPmij2OSB9WdFxWvdGhC/hgHA
ge+hq1pC9bVb65chO1YjRRd2txNl/eLCte2pAUpTu6a7VyG//qm8lGfn+cI2uTkH
lLUatS0UJ24Hz+KGOH46Ahu0eXAV59Id1Y3GCpnJk6EixF3N2vNhJh0IYod6pLQi
A64Wc79TJbzwQpQ0tCfnQGBCzUYs55GBc/9JI0loXGJPizcUMl3P/EYiFM8NxUfu
CzfSXCOH1FjOwK5NsnaJ5lNNXEaY5RBS3hNqzPPj8QluGFCD8MP7mKVpeOcjzq23
QKmXFvKKjExuOu64Y+WdNewpdN2EKGtxtWe/xPZI+H337UNfw+YZ5gxpt5rddHJd
juwASQlkdgz8mJCHpu7DwKpOqIgnSanQgRqzBEDGvfeCK6y2mFwso6paaXFNEtCv
CSgW689D/ZSKX9NbBfEEJogKieE+mmji8YqEQcuHLfb1GqMS1dGEtpMx7lSJqvks
c7KWuCIf4ZL4HZLFHh1fys+mzngPT2ukLrpLMOqlJ2BS7FacKHClHGVgEgwkmxzu
b9nrspEKllpxGIM5kpMD+U+HFUig9luJh37D5xpe+TVk7uwhAiLiZ8eA8rbPbyjD
B44NDm8oQRqTSl/yHlVB5dLggwvMPZf+6+wNgzCqpqEWdcj08yWalM294K0zwzCN
P/1WbuEDsykkL0grpjRJ5BTfVeFzvgomgsj2tY4p2mirlCu2lKEsXLsFHWoXShfX
++LoG35TfGdJFDUkMd+6CKS9NC1alOQB3Q6XxP8QBHqitQ4eDdd/SiDhNE5UqHQK
u2rb5YHb4Nv4WIeaQ/G6akGJG/j1B9gIYoWwOtRPwvGz56bFl5hK7s+invEOjXvv
DyZifzSLgzy8NoWucEan1X+OprdyWzt+U9i9UpPczSDkXWnPPRONXld3iUu8nAfD
RAoXhEdZnECdCC6KiXy3/OPfVjgwbw0tHBO2oV17Hq+lPetr+XZLlwuJpPlcXpVU
k/+D2ODwBgEtcXLj7/Rx1nABTxn7Vvu95XwYre5XkL1HzSd9rxQPL1eA9FV78ERk
KqtgBv8Ro/JyGdBQ8/KpJdpSod1MnNEc61wUIeO+VI+HEjGM7W2LV7lixSAFVPPg
ixeTqqPzc31MgB2Ziz9h/VumSZXBT2j+VxWvovxtxF9HxAEEgYdePSvAo+Yk5RIe
zd93TZQeAxZ/G0+TG+yUisErJXWZ6Ki09J7Z9PNHNRBpkwtUukcCfRDlzaNsTCU7
N8XFsixf0wLtY8Z0A1JICBqGIvLFMQCU6fGZSxfLzpJuwarA49/sjDoFpxRU5+Ir
krRzIUwmqh/AYEssBQTv5070z30a9V58nvxbQNXwL8DwqJJ3HFVxDNjzWvcNwhMD
JQgV2wmtg/IdJ0iQYCBmBnevsMzTT8vHYiZTHavkwIJDdbE3XuI1UiNfKgApZqna
XBthWuXGD4AI5SvXoly/gU5KeFXMbE9USI0ecudbY8N0XN94k7fp071/Qxb29Eic
oo0aI5ldkqXyXDqd2hNMwh1Z7r1YSAACwv+vaH5Df6XfnCJ+r4g5NSC4s0gAGWsu
gd5DD/+4VRgsuf3ZB7C3P4n2mz8juW/zTbBI3RvtnUorIdKoZU9CzxpbNmo4Uenh
51PPiYhmQ24cnXG/vac5qqZNAyAKruz9jM58A1JwI5hNmsuQ+oy8Q0mJc2VCrPgh
HHSxKfztn4LDKQ0JiJzNc4+ViQkr4bRfWOTavgmu6REcy7Xi3brSlGsnG8POV3RD
iFtzkwM7H77cX2EpTtMbseiGfeYZiw6hsjTYfkJ6JYP23oiPQ0IYuB/xREfkNu9M
S4FQYLY3DU38Pn3SkU139WOyxuVtGYWDtofHRJOobQH8UzOmSUn7/SfRgPbsnNnI
IYpr38Vo2RnNQI6ddb9Dy55cxgPQ7cCEvz7Ef8h5jIkuoIaS9gaa+UBF4bEttux3
OFfjmL0KQlOgMCov+VufjaACdZZPySWICN5VHRvQF70h8KbUCVwCLK1D+qeGaCcN
Z01xicHcvEV78NhoPjwjcA1bgMAgy3cN2Ji+q5RUtETDHPH4LHMavg5epRFWC9d2
9iLEKysVQHG5JIgZfdIy3mgKfn1XNg1ZQbWS9TRTRDHWYyInu5YRLb8pLK0wX5gP
inHW4xehik/tvyP+v/kplw4vuqGOUJQy3EVhE4qwBJqlhsYWSTJ00w7lgQaFWAFc
tQRGVv3fJ1YT0k0BsorBz/LvMC8bufBscosDJ9sbg48o5x2Ub9K+7tprhVkSFA0y
bOrU8qz0O0Xh5UwYm91FJBjYMyioN3fBXHFAdPXqNmtmXwQSoykhNxpVkCwlvf6S
zav0n0m4BzobflfH6jwvqrbF/x5VzqUzJN6P6Fs6a2sTJC31ciGxerb6qegncYy9
bsdAtMIO1ajIVcOiHK8e95/LAem1rMQtGKeQHiokTJAWkMVtfeuvtGo3bpCLy+7s
IEd0dkEhJQnBf1OfbYzy6uFfD0W/1JxI86I4tmQVHLkTSumOBxKVxzH7BhSSPF4R
NKyQCqoUXXu7bP3kXS+EapkFh6LwftlU0xrFsqSHiGvjQVzGaAojS1wNR9PjUOJu
VfJGMDVQodVN1DZ1552H5QewzRZq/jjinXDlTIrxpD0KN1er75rrJsvoSjgblDeY
+YnjGR/ILTmV6VFRH/9pmcFsfkAzhSjoWaIIrznKsfMl3zt4c8Ln891RiWLLXvee
Jy39ZvMKd8v3hH9fczLrCDak0cjD8EWqxbYROX4nOmY6tK4TNpqxif4cs77CIZuV
RpwA67FCalS7+LiC0xodi+YHvBtORa8w02E2t+FyfrozB/oADSggDNPHx2W/WZ84
VPcD9Ilbe5g+2HD1PAG9feXS4xTolVjUJ1rQS5xd8XuAK1XXk9XhjDMuZlhl7e1l
/jQIBb5klqsw9LBYDah3Wd8ywjGbukwYIzzNeONtFw56vzw9249SaoKY4Xz2pIgx
PX3sOFbPQdSzekZ2q6JaEPO4py8MHG5ZuSVYa/L1hTYrOnMB8FYwsNPuCyqmyzlL
P1khDXJFaKGgT2nqpxbgufcfByueaa/zLPmkyhLUVnnRLQD1NNgNf4LUeW2Ryk9+
lIP514bx/Ebl7sa3QnQBLD7QlvjQG7nOEBq7gpwMYN2hR/afhWyNoI7XtO2gRMXw
E3Ocl0okrRd38RqVnDIz0jQG/rN2ibLgstlga3M2weLWGjfOGodfxqofdPQpx991
077rdi8idRrSVEHwAVIPHtIEmc49UP2azl6gWaGiiXpLLY0qhUTEwDssNu9ifgtb
X7p2320kjuhc/n9UEZoNp6lvhnO0Exe4lgjNo+xg7+gJVZy6ksIkZ3hawuf8bC9A
vCnlqvV4aCEF/IpiOsOplmjcUOxvH8X45cfAigUG3L29/qu6/vJBE0bzLVHVbJpZ
/MEPANCuXPNzNPuuxPceFK/xAmWdHM0cbD6E28oJIYQstbJJn/9Zuf3iyNMCI+j5
8mXkf41y2uKnVdh6TPAmqWmobBlKVDpG5zFFOudHSx1IlODf+SkR+LEEWipUqU0c
zjEnymJSsKvuKp441eeKB/6bd688voDdCZfFRALbx59pFQfwT9t0xVA66Xd7HlAB
mEOQ2szGBqDmDIuqCuNE484hFIRuTupeH3g7B5FT8oSzgTK5WSEkhNldLZ48HVic
bIq6H+IEyXmmf2Fhvz9iF/OZ/I2M/dJLk/25JrHC/zsDNTUKCfDWOHT7Ys+WJgmI
NmWtgLXiRWjyjEPAxFgXh6bcl/R9RBJSvy4JOJPpquDmdFT5iwleBOEcoKucVWXo
dOEz+OU906HYdvAk8dIddsDFC7ORJlT/chehzeUnGeBHQDAFSpzxdXtKKX8amKeZ
oi5/n3SMbj0zpXaacoGboJabLrETuBiGiNGmKKyZhCXP1WxtJSbxpDIVsoYjTWCp
tHutRCOKWDdrSDDHiaznyRH0ih7vp0u0sTUuA4av1hn6w4IhrnGbSnilkVNiQbtt
PFndtvrRVaVVi6KY8BfPHpEvEli5b3yjDdE1iJGuCGdT3bC3B2SrlzDn8YHqK0PX
yH5eEnSDcuKlMYFgHpMex4vmUnJNjl2AV3XnM+yUxnGnbol6YbbEkyXgDv074qnZ
rRonm3GFuDmcnU5NJCmQTtc3OckMbfJ0Xfgm+r10xfSTDjMSiHRKAy5RI95mt7TN
V7S0jnTd7+A0Z8fuFOq8qvy+tmBjd8vbkuUneqiCg+and5DVMJxEm53B6FoqOKvC
hpcAyXMFzPko6tdkuIypsVgtrNhoqZ1pLyXb1kw9XXthbCokqG5vQHPX0Z/xT21G
Xf/Ih6nBzesvohj/uU5I3k3MZtdYkXeTlQTNQih0bjFjQ/HvgAnDLOfTmVuRSnu7
mBsPQV8AN4WV+wc20KczIjBevI8AAgU6Or0zwZPRh5OM285yHx9Hzw69KZpyU6Ep
ODwJn5Tv9LLKCVnQUwemBhjc6XBuuNNmEejzvf2KTyST7gZEa55zJ7hbHRN3wjUU
XiEzvAeVfIpCWSiD+85vzcsSI+TH0ZbNBnAs+iffruaelIf/wb3iCYX8svqYMztB
1F01L1lOWasG28imjSv8uaJ8rpLRYnzZLowbsQM4wdzYClaxSB0GVm8D8yVfW8wE
VuTu5MRhndgSi0e2aPZilOHoxHctZA96hmEJYaWLuip+ob0zc721qu3bWqFTCje0
xBTV7NXCRCFPUQulmUVaWPa5xkKspZqdYAiv4NEjHz8Q/MPPCC+7eYZ04nxfpcAF
HKXHFkBbKxBEikW/6pkKpyJdVt8jIOMpdeEz78H0eWurLQ+XYJcIPUYRCwCq5su+
IRauTcUe68TZJadEpH2TjPFqc7qjuzMOVcrMQMJNSUE1ii2WKthW0fleBMbJCMOp
IxHqcyV0Q2pM3Wz+g/QkVljRkJ5QNJUynr6hCr9ogA87MmPMvdPxIH7nMf5xyZnL
WVowmZMbfKaFf9KPj4sb1STI2N4hc12ILfDtZXNvDqG2VHFjjZYYJgYO0g+VzzIt
buU841LgcW0dqfmB5v/WlSq7jjhs1FOvPWJswgFQ5p/OUwstcpFPC5uJx36LxEn6
WKheb0XvDkSUJxiXgXBVJH5xX9WkEzJM5DGMw8taTJqnZAVXciTjSFfYN0IEluvw
X+bdCRN5RV3l/ur/gMK2ZB2uQ9s06R10YEQ0vc9kyHRfY+Jo/XWLp6rFmYY+haeH
/waSaxOEiFhUVYG1jPTyThdjtrtuMyhy85nvQkYSI7u0G41Zxen7VTXfNCAX6rhR
IhjMyJgTfVxyhO+jAnpEnsl76qcEw/2z1VKXQKYl88I/xjAwskcZYHp7pIiUrWza
TtlIrnSAtwau1tyBH6OdP9k1XUzEjZyVDLzumYCzDHgzCtiBLC4pKgwsff5wOfAi
IUQuJmcDRlL5ng8w49oOTOm/S5q9sj0w6ANNPZ7mSGkAdKH4AFq3ubZRp2WNkjet
Ycv7pMeChn3NKvcNe/0JUCRJxjHIui/uVOylN7x4BVLF2YaoRIuw3DW1+bmHqkLA
8ubkke+TDe7eC3cv3Xp1M4Fa8dEOsFINv4JThjQrDtk0I/mgPs30eWB1NGqAeP/L
KyOV4nDP8NPvexEa83o6lP6N9X/aNG2GMfS8G0ZQB0nW3LkTNpaNyvaBgUojmvGY
oH2Jg4k07QntZa0mxinFCl1q/U1xBuAMhNzseO8ivKvwSZyu/M26VNtXgi3851Ds
LLlElkCz0KSjolD+PoZJBdlI0eO7v6EKIY+NaDW2CmVoPtEpHW/V17bN0YN6WI6M
PiLqWVlT6ll0hT4uI6a+qJcqkTCuzmACke4GVZiGJdObbIfBegFhrUJ7ue0Aokcg
UZckS0KE/w4hMpSg8pkaw2p7JRjow4dvwMvzbu8qiysF8ZrM2MPonCkvwz7eZf2z
z47gVR6GDfEVcbIkXTLObndUsWMrakze9lNa1Kr26CWvjukQoWzMlVn7vEYf/1ca
qg45skFArdrw4y622gtwPR7HrNQ4N/N2NBgv9RUKgGApp7Yx8SkHiKnF8d8YCiEx
1cZNZXsu1z+WrAddQB9Hcglft90q2qrpMg1x2F83vo62Rk2zimbknrPECumwQAdA
E4MR+hgrNYQ6YYg7g9+YCA5c/zqoO8bpULvdXUmvVesQdmYyXrQIfi17gh+A3VsZ
yFLGPWjyf9BSkP00LBV5egtKwDHvL/aQKLK+pTCColMkozJR00lstwsGF078ctj6
z62By6DhKkyqAsAiPQ0/Kin3WJv/bjnYQpgbaKfNA7ASi2+vT2Z0v4VobnjXHIle
CPEFjR3HK+HPC8puxHMr095ACbHRz5KkvuH5ZOz892GN7693z12m5aY7VxFpqfNM
n/4TSvlkptxGsCHMrKfjcAAVi+v/4130kpHW6jMZxeB2Qb0SznV3SAGkdnrl7j92
MlW+HuhKOLBkgZEpYCinVAZTiM4RW5ODNqlLnJ8hZWe5S6vHjAix8ZQKHwh6Q3kg
u1O+P6G3a2Xo+3mOZxm1Z5MyCaxlqAT94WY9X2j4cZdKq8htMLm6YJGC7MtJ8Vu+
pwv6E9QAs4GO/aDyDo8GRiHD+K6fpPOu8qrDHOShKRfSKb7OGem1pNpmgj+YbcGU
h9D+XZ9XXqRA8jsC4ePh5gcJ6bSHELYdz+1rPyiMa3H6Bdt1melDFy5gzH1cidtz
zL0LNNObGe2z6JtJzG6wDY+nv/mRxACFhCSwEqqTfftu+ticNxHnyIfp/SmOdYNn
/TpXmRfzGjkPsjqE0I+mxxcW+uoKumDTSWzj2VaP9VOSBkJaxlrus4l4YFiMWQgg
VgPQoiaKyLyCMZbDfF5ZcPjAhF8RyDOVkZ+TGwbwf3SvJ9v2BP1GrKWzOXAzsqVq
fqRU4cYPL2n07qkgk10BdYLzJquMdM0g7pzySjyNwid6Cs/Aum9RCmNsD9OVWPS3
IPuiI0qK9dvIz8YJYsbn7MRXR5BVIGRDlT2JuVVUthf8FwYHycoS9n7Zigy49Glo
YtPGE9VsJd5UahAxBGoxTmjdadHL24V88LV/TfPy0WjKDEgbg27iMlqzvt9vy46i
CtU7IMEgVAYZMF4tvhYf0ww3B8uXFkZ+mkuqgyF/gcLyuMwnxXsElbFRLahA0RUS
I4VVXFCEqqwB9CaIFuspdOF68PID3IfDAjmEbdTx17xRYR2szIND3gqf2eUmmtke
qwFjuhT+RmujXe3vmjzK6M/cMUHbIK2CaRMbj8jY/Oyjqf43yeCsV2cNoJEprXSZ
Cj3IUrKBJObWottrVY8jjUS/5ZZbwcjp7gM7KWknfnL6imBfpbfhhgaVog3HzNZL
8UUuVMzpXiVIBDp4vPWvEF/RxgVT5KJLEk1+utfVDNnVMwfQ/i8VENqOEqUtBYxn
okHWjVRnq5lU9MSTKRui1IhxtNwLspF/DzVodTnA5ijRgU+m4z8q32kUDVpWc0Vn
FoXe4cj7dTKmrNo89oQwcmTrvvhrb5qUleja87ZrI4ANlS3Vj5iLRZf8KXzyMoLR
jGypHFuFf00jAVrvKiH9OBBFcpEl/ZMg3BF28Th6m4jeivPPWvVwnHlEmwFPyxNF
721TdJ31a+6chBX2g5A0/9gmXfe6yCY9c1JyDHmi4ftB+Bz+v2/rr34ywpEPaHVG
acf6g44Z2DuLMOmM8NDasymOtqnWKDJRYT2CTR5IuP6HNa5nbUSlIgcc1Rre5LM0
3GdciOChGHFEFtFmBLl+hrV9xdEmEQWlcIVQKyK4q1gIxt3lJh8K0OoIKpzob4Mq
IlMKAu654GOuAnW1YaqgKu7iOPyrMouNXYj3NgnlSd3TR1efDgA+N8zNft1JHwJR
+LpyB3DAskmctiNbNRjyzrZI0fNWoUnoRY2YJHeqKKmIDaXe4cmXGnrFRT1rWj/q
OETnIEB5HFcNeNWCwIE0gD/A142taqnETB63Ke0ZrKYM6DanLzblN06NNi6hiNKx
qb8Mi+0C5K8ypIhgR7BZhlmnjOsNr/8suNZ5wTodmgN/jCf2JqH0R3owUmGZjWQF
2mfAK1e7xvNwjQod+mtqmXjHDX41o0vbyvIRLW/KhyRyv9suYy27L2X3k3G5IjeR
pSOF7yCGFmMoczjwZFNq7xTuFom5Gs+eda850CVlNKTFzWpSc2NLup7uR3jD4/Rx
hQXK+LcvcPMlDCDmP2YbQke2NjDdeCaq+t9VwjwzsZ4KVFXL1epSpz8QAi3HjOWG
w0TXqtTbYUE/gdNkzejjJRQIsPw0yPUNht74Et7cQAicNUKB1zIHP6E4O8kRRSQk
AaRPP5PP2IEb0mgYoxubPOP1oGXGdlv1CfEim+dK6DUGQL03OVuu6ptL8fr7OXDJ
gy2OYJcLYsLXT8RX2lz3y7m1xr6QYXtdRheq+Wz7bv+7EWbf2+H9UdfZ2Z2Zegie
hibIl8BOO/tyFWw4dSZrQQrHm9uW9tX4A52v614NV8iz9jazBSZDjEnFDryvNRUh
mCzsXWuZRzSPY2TA37tnTsvggj/3zOxsEmS9LfC9ZbNI0BztU4r9DAUkm6QhupZK
QycYV3l1EZIJa6H+NMShOevwwIKAIRqofDSHLnNZe9rqcOJ21nrjyiDZ29aKWmo3
j0GXbxlxhb1vduA+9dt1FlqRJr55/Pi2N02rH6Skpaai3bRhKwxlrUhupEEVSHYM
73859py53hFNt2GB+2437LyX+U3mJTJe0lEo3nq7WR4TuNHCyETpdWko7yBVOTbx
gK+/fNVLWaw6qjnStqEg3VKr2XlnzSUpSIVk85hSLtD0Cx4ri22M92BndMX24+GV
iLxz7mWAMHZ6O8fUxPGu9JLMbDE7DSF2Hlu7D9z6Sn5q4XAN/ItLcsKvjIXI57Ul
Clpg5L3/vtLSrhxJYsEW5+hcRa6r6vzEoKXX/ezX5He/L8CgSE6eNXjjjHWwxbKb
bcaZBFsgiJnhtHALkmbf6tym7HwkMbJBKJEouNTOH4QeAz8zTIhkSbU1brApLx+q
BDNEL6ZB06CeIWouJ3TCzDH2pwYHBI9AFTMKRtyrfD8FkIcKolxNGSWLKlYTBKYK
OGbFt6PEB7saexXzFadwYfu1xXlyenkHIx4mjrGEUZg9z4fWqvQZP7gL4nQAzY0E
TbS9xoHgO94m3U/0hgK2QR4iY5GlG8fbZC3xX9tOQ06UIaOfVa1+6aAvewPbKjHz
aDHR3k+NbkhSEfenxp+creXhN+mgrWwD2h193ALK29lI3an/vlvAV2mKcRDFs9qt
1xmmWKBm9b0mAVLEEdKOvvT4JTzcp12bs91cISASOdgmxKM6lvT9juLSlxDgUDwT
sxaiyT21vDMEtwfoq1KDhYZujX3QPrXuTe/VL72rCRlBuqSz8d6lBoQImD0XxhAA
VkqgrcwBgBDbbC21qTqkoXwlRPe+3CsSAaOT3geQogLzrnjG2H1sFhr/wfqittGm
uZOligWwoFEB39I7TbojsaweItuKUUJ8QfIe2p9Z6DFI0DCNCjhDzHqTKElp7kYG
OoWqhYfrHEFmnoifqGMmiwiHrmGCl7B7zZ6iMIcH+wLud0qUPHWPhwD54xubKyrj
kb8AlbMFGg2+O1A1cmcfDKQWfcg6qcB3TL6E47JINyp2+QmxWvmiMd74c8XzS5Di
qMLj87/tx78BJjz00Al1IKn9Dn7NWaJxdNdBmlOyLzZB3jSSDc3RJwteTsNPaocd
waQrlH++ukyxpGl3arPL6Hb5wLkyWxxo12p8t4+k9PnT/ouPCLwDUSQI/LgIBTci
sacEgKDn62oHvBtE42M7LR6GiknAj5nqsBYjC3UKQ/J4EzUbdkgxV4Arn1dSmF7Z
/Z7XwJ/OqCBDHKRPJR+sN/14neQXzUS6u7CFgj561T2+bD2TBwWnsODjowxyQkLR
Ztc2/OGz7xfE6K6TBB3t3+vujBrUKs/fbOPkxJWlltkpQeY2KCE/IQAIcqEx2v6q
CXvANjstu7JpNijsJ0LO7viLkFuw7MO2Cww4qVULkmv4NatrLtzW8Lmb6L01JW4J
AZCVsZzQtcDiXxf9tfWtmKbL8dbADHRdkYqkQUDh4QvIegOjUNlaSr9FnQVQJglo
sWRuCtpomRJSe6wInh96QOmCdaZZzf7tWTPyRI1+Hm9leAU177wUvz1hgG/h2mEX
pZc1/EZrfkrkq/JeZrfJqq2r/nIeRrGH4Js0Z2CH4p75NkCUzjR0mOEPwf0yFk/a
3OaelTxNHDyTjruiqDEt4RaD4xcLv7LMali2s4RscZFwy1y75IRohYbBc1cPiAbj
915VQg81drjoR/9bJObxXIKocUlQk8UnrgyLuW1zOydfG+GteyEsem+EqNnLULxW
WruRD+2/MyO8dbT2JjEKCnkz8IHN4Xe9y96dsuBsDtIEg4RuXzqTXIG+6JjXgtAT
aY4QRKyVUWxkDOYDW+RiJmAdPzuy9uyicaOUrBxgLH0N0IzJr/ZnBRu7nwQM3P/g
pxMwSGRHuEeLbTqJtNif7SY6HDC/+848JbcaiDU3lIn1bEWWrR2KLnFVP6kNxdCd
xkDyyGjamSBz/e6LluddL7W6ViWZnC6igGcR0STLGLQNCeDjtc7KbKsPl54Rh/te
YHdb5CviKKMv/bUsSv8qhmU95wxfN6RxwupoJgnh051yg1N2MkPP5/y4ZdOJ8GMD
LXEvlnEMjzELwtKgYhz5T1XxeF2GDYAGn1wY39HwsYefKw0zDn4MtX/DhPUO8VZK
72F4j2AsjGzy5I97kSnlN8ed5cbUJp2oJQ49Vcnt6hL6KjSV2sbgw5r5CYzqpOyt
RltfTHpa15d4tQKgbgd4yKw71XvEWUk8ccEmNELkVAqvL6JjQEhAPLxGKkqF7eyT
xSKxyM3pWFHEtItdCK3OtCaIo1tiTw7UYzUg3IWhpjwRHddKEBa7JYtyjjThRjo0
yC7Ad9rjLSSyXuknw4ztoPmBTgKTuk/IUNsyz18Dj95nIfPCLjrHDSo1PNFCoqMX
ipTH+PWo7PT4U3oQqHOXfKhEoFmJbq2jzgYWOlgu61G/gZtGY4G7rbG2shKhdpG8
ogbgqPE65YlwvN2lVrCKQQAGOFMEDeVdnYVt41OoiSTgxHwwVLDMoPcPsunNMpLq
OnWhYhclO4aOW9yzm8CvSGoFna1bckDP7DYjx800/esibieV+mkWbmwva1Hfn6M8
Y/okOXYbuSzKEQgezMhS1EpgBTmUEHOnYXlOJotRTXFY5Wuzr1v8eYAMkIyWfcpo
nyjnFai8OMfCXyf7Np9Z0XvfF5HHl0Au1cStUE9u7QYYPQsI0VYDPJoXeDfwifzq
s11UA/70fnIZAMzF9dHfson8LO5KOVP7W6fOr8j3GlcpqXVf5krJguFEFVR072Zl
vzI+N0rwXMJkFDNJZw27ybjYVELvA17O+qXetZ3pja4BxR0Nz8G98fXMOUp27yut
L99rsIXtNjhmBVzsMDKyALhrq2vOfYEDt8ZftBBmxEtdI+//Jo/4H+e38tGz8cq3
2jlOMfOGb5Y7ily3aQgiW68jaMnxK+EYk3RiX7+suMdgChP467rgnzN+hYCR4xB9
FX1vcSmIXRuYCbNCQ9uEp2wU1qopCN4c+6YNQJ7+htoxhgtjFQGonj7L6WuRVNxx
k76WdiFn6qMOYoEEGvNzoGrHIsNf8gsQ5fAR8ALEpW7nd57obHlS93U5dPqF/kxq
RUXzCw8ZA0og0kNeheslgkoUrQmRTd5Bgfrn0bB/jz3MiYIxEuoePwusnwVTdk2W
498djKLhavcyPeh0Y9XTAEbfdql+pvnDgRKKamqnO33tSXOLSjH2+rX3AwKGewrt
l4fLzNTBzbHH0BYognRsj+vdaJoxhJsYBspuplmHxSCF5Qwv0VXSA993A5lAEaTh
ygfW8irtE0/Gwq8Q0bVw/ZwSUoPqhejPIx39Cpi06Cmn3v1atPBV9d3M6FwYKx6a
yeNde3i2aTBHWP8uC/vyz28BBsDw7yQrNNPC5OFS8ZKywDSZpItBPF/Hj50a+F3f
IZEdxkF3JEejUjPzciXPORQKiXC1UTDWA+GES7NPI1KsgYQLTfRYFBMLpyQ0EaTT
r3Ed8iyFI2znvOC/40BP4t6CkXutP8nlHFFoYKTgN5H2NkYqZRhFkwanrO22+1y+
HamkR51n5SeXgYQZICLpkwYp098FfxU3f1+qP5lyWCrogwELBByMo1RHRutGXWC1
DmfYZ9/fmsVBIOyKrGlVd1yI5U5HRVLexu0gUOVQCXB/cE9TWAZacgsTnTGvXpJG
ZIWDzublzdFCj+cTARrhUROJhdHmW9h3XZWqHaw7tyFu3+9akERu+2uWraH2xL46
U3Uv7QcaRLBTUvDGGwxvJe+k585wyBC8VfPyDbwt0o5+5hmektQ1fVvhq4vTvlR/
O1wRebzQPfwToQS0NFF1ZVIEB22PLNn3J1oHJ4zYpE9L0qnt033QrpQZXMbwKqyZ
pMvYcEhnF1x8vFDljysTkQl37BAn7YWFJxFrGtJXvU5T9eIRnHwDMa6IGjQH5m+V
0988prlRnynjtg4H+ytkH7b6k1or/TJlhrZKL1DrGu9KY287uCyqYCXoexLswnP4
feqRkCP1iwsbFIJjJYN4MHKcdPCkSOdGRsbtUuN8tPSan5EfIwHwY71pMSiLeDxK
ThCOnl4khM4QQ/buNP8x7yvX9yncdy2NNHnKHbisFNoCVpHa4TSpxTs0NPADD2ln
a+HZb2QSCyaJwkdzb+Z0f7cwv8DNvYid16uQZNdVoJ4IGgvMYvDZCsf+bEBnfLb5
DYnQuDEO4bUBdt+zo+KNPzl4Z1ubUctQ3bV7cHmMiqp/WAwj2QOVZ7EUa+gUcb16
sgK032HFwNP/VBJKhco51Dn4UsYkMCwCuF1k3e+vaPGHx6bs9BJ3YEqW5Y64hU59
gTvXBGLUf1Rtk9/xuBizpA4vST5Jez7DnYveiARsucHQL4LAK3Ul71oNdtr41gSz
3oTVALjBwgQFJ0FVW9Qn7zaPTRIjvRi/4S1ZtgjE9/jPa20wOpl/Gm3od9yv0tpe
brfAgBZEBZ2gZZSlyRH+u6HVhhsUNyTlvl2V00KdxxKzZXTR0W5g9rX1odJSYYsN
BLKWIbe6hU+yt3cd23ZAFAjZ9/fsFcNpS5LzGGMCQqdGgJOm+dm0TE765z5ruZ6V
cFkgQQ2Q33hGDIHeHIfaKr3S9GkZdgUUmYZ9Eouf2cintDaoCNq4/VUSSiNE9cPG
zNVN63GpbYlPIt4JPhkuA+VFeBCO4GmBaaXZBv8576WcSOzisQ+QEekSdZt8GzVz
/wd1847slecx8/mC59RjgsrfCmGNgpATXQPMH74+BwB91apLRMC1J76a5GafiDKi
WG3760zLiyVgPQYlmjGl1u4eZmOHCUNQLpUgZDwJJ2dpX3wbh1ZaPy1qz1OjVySa
84z+n466ZPQod1X4Cw5osumiICIbdMM53VNm2fESgcQP9G1bWQqBW41N9b6AWmoJ
dBoEszHM6pcGjOFiVT5T4QB/Lp6ItalvEK6Nc+Kt7kveNOuQpUV3bOZ+w3ClOV6Q
5JYLvJwb49a6D9eccy29ONqKJRRb+cVnRKgvxpyEe6tNhXCK5eRfWJjyQqZCvrzP
rWDd5MaD57356ZM9qSIVY/OhcClBB5zePI0m1zlCIo3q++gmxdOmhnNuKRLTSK1o
zlFo/jubBG+f7gJ53HB2XkOnFmJQj2we3bF/P2fc0rWPYE8bJb2G8SAVQUyqCar5
L2EiyEk/z3rTQsZ6HBIIrR7wmvpIPspw1HPyXzvLzGlJbz44CmWCieRClvMgTFSZ
j22Jr1au60iti+jFp60dk13jK1Q7KzK91OZTg1t1ruYNoZcKT0W2SDxlMJuIVHJW
HQcmWLYLZbJ/UFZ+4rSyYHIE9ed11i6O9awYepVMhvhbB1vxkLXpv30Q1VhhL4n9
0AXn80HKZO3/cZ6BHWK6hUeQLlve7Fh+VfsN5O7gezF2BQyRX3l5A06qmU3cG+No
SaKKgO2o8CzA8I6c/Sla94Ab7TzLa5Igv5qrhtEr5Imdhpl9cJhsrlJe7sCSTEOJ
Hti3nVyuDyYDsFFcHiEpsW88COuTEHoQ2D0I4GFmSiURPc0XvL2v5aq395nzpH1Q
uMfkUT1uOqJCB7pAk6jMbq0obGSRmIvrcqY1w+yT+LxNCZIR9PdH/Lw6ny/vI+Qd
BWwZeZQqEVgbifJUCL583E8LWY+0CMnjNdFq7YX/K0R7Bo2oC63CWJxj7t5zF346
bt+JNhX8RaWeUvMiB95/jyNqsDZpv4BELbyb7pGMIuDNTKdvnnCw6TbraEJZHzEf
RFxo/avtJGoyVHxIUWg45S+2b7NdXAjFB/vNiqcnux9l8eiw27GhOyLFFrzUL6Cm
WOr5T6SChmHau41soKFMK43XByKPfMKFs9/TB4+ePprRC9zVKGbnqERgGj9S37cm
/niE22BDAmsdIzzcAppUWvVmIMHmTlmNQS4gWHgj8Nagj9r980IjCFW587/0Agmw
GUfmZjhlTa1rO0pXp95NQ+cHTvjrc5e4KC9QZT4GZOsSZ15A8uYZTaIIwRkimKaz
M7LX3zWmQ4vll9AxZng4OeqD3l+zJuT8a+ROOqO7UJETUOsr0qVgpnQKGrWIFPou
AZKv4KwxUQZdoJfWf8ujk76vWoGIKBZAuHC6mHmfSHf9ffPLr4oXcoGXF1j50YIs
RaRrpTpQTXfNPPu0YTSXIffoXE7Tim/cGIjHmjKVkHwiG/hHv7fyNKgYggzUz0SC
uNzeaDnmSRYeVSZvmC41trJwihfWe38ZwsQDV3K1QH8ZxQQxtfi46XJVZelDnZ6A
APhLqYi4q9AeLES7BX12MAVNqa42g6K/SbZ/ojTCXRjDt+lDDDVf/IVi+0IPR4jT
IvfJRikqZEETKnVELXPdaOjWC31QpP0eF2PpPAwpn+IFG44BMUmcXFkArSNNeGGq
46W8UDzqGsn+hfBxuKMuKem1mTAX5WYw2ekw4fYohstkaNjPCL4grMtAB8whuSaX
B3JSz44Pj01ZfjXYkqNH8qdYvqKDAFx8+Q5rftgsSAozaVPYR6cCGwLKFc0wqQ80
OK4rChS8mXSWQ+CqickkRxtcLxWyg8CmimILLRBAocOpyl6qHzlxtK5R+OCCLpBG
p5cIOObi1AylBlA0i2kr4FlQKYw6dsektstYZF2/w881VLY3GAmfYWVxsmnWiKch
7V5Pbf6Bz9YkSWmvD8xIas9aN4nPSK38QQEFRlhTXcnjczuVGIHhBj7Bna8qm2Wa
tOdakR2EKK1LyiDSMqEQNoMGTi5Icf6WqFlDMc5fygL0yBzg8XXm+MInqdYmP98t
J5gnhTIr3IyaRmFsLd79SWWSND+LK+X/Iwv8r/jJXDfNDtiv/we9T5lOgbN3NWSa
C375y+sLFBupqgSXsiRMHpjqVzV7vs7usx/FyugZojtlCfDhjGcRioYuUIwrGcbB
gVrMHaCb53QEeEGeJyKOBHvgdCppXXXoE7RJn6PqhHsU/Ard1pTuRyv3nO0mjdK/
qi/G4KXbjAE6gCmJBu36izaKrPDHNLW79FuMpIl/IVU9MhlqHKRy/mgAtnXqPAq0
o2mnMQ72c9uVaJYE2fe5gZuJ3fkGf/tVPmZ735GszfArlMcHWMI1pZ0AW4DkBZFo
C8HLvLb5qgkGZRAQMaXqL9l2agB0BR9AYZO7pTaRcu2QVCaTls5lYmrUn7q6rZcn
2oAjJDGaFVdAZo1HSaQ8YYskA9NQ2VUg+nvYVd0tTE967fdzxwpmG1nhKrRQJSEy
ucbcmOKc0OCp9zE5KgQlyW3UwTN7GmLXIz95/wWG/WvMrDTP3wrScvYJubtr5zYS
ZwxhJF9An/zsmP2rdvRvm3kDTPke2/euhwwJR1OOLS8xyc48dLFkJxVtsNN1P9l7
DWdCBZUE2GPq+3WQiH2ZCogo0lSFlX9MSsrr1zjDxsYRaabQmVmhYVv9lSxRnR1j
qEfv2f610Sj5BFYBoHTAvlpmmTetJofzP2Ur986zT8V9KJszkLzXJVI+tt5PsgPh
TtZkhS0G9EeBpBFGPvyImTapKeKxcGiwXaUlYabiLll70W0/l/W9KXkMhy3cYn6U
HYO4K/FyNMocKljT8CYG0yOpVX4YbQRZPBMtG/jYYJ9aoN0AohNK5SiEd8kZnlLO
W3r3ViLf9F7nG2Rm6Q9RmC9sgNEd/xhEBQOEcf0qa+OgNVrTwzqcdEvBNAYXI20S
MJJY4fNcGGSpvYPix4K5ay2rAuwLDHLH8cYeRV1IrEL+wsMehORwGnN5pUTGkD3l
TSCOjHFYxSuu5VM+tTybFr4SDfYpJ4THBuroGlkvQmTGqOweWf+S1+MO5PDSWD8u
A7I7LdiaRxvHtMs9PTXHGKjrtGPZU4FmoqdkZZnfHrMnp8jZJh9MGYclUUFwR6eI
fVBkHkVomk5D15zfAsrqXHnTl4jlAPgT0+eT3+51KRV4Km930Tfk0FOaaQKI+KDb
z5eXHrjMwhpY39y1trwn1v7wrH1goWxtn6EKpl4tH8T+pvDD2yaeTX3pfdhhidJl
kU8J+s0OvxAgbu2CLeaLWuBwpY5E0ckwIjrSvI04Zw3YS/xyj57sq1MpU5o/ggVl
epnq9bze23WDrHpoCEJWD3j4zCkn0oyXLC621TR47QOOMQK1fLq+xartdRNLwQWf
ZZ2cCAt3ffeSbQL7NeAW8cIZckb8w5DGsTKubt2E/uyKITRlgktPLHf8mzHprEZO
wPzMg32l+2aKTIWrJoE8ChPl9DB53cfBU21Ze4zrCgwV7aCjtxQC83vXyBUAqK9o
+SzXdWOtShb4ZohyXTtlzkMBQ4tJ5l4VXShvDudj0KICF/0PQO4l2pNIBfYvfUZ8
rRfvetVzYAg3yx9Zlwo4++TR240xsmedFxea8FErDSL/I8R73JladdMA8bdTFsxy
Tgtnu3NVHL+uxkzijkzykfy/uzJI0zoUYtxndcKPx+hCi/j8iv+5b1ciTSir6csF
DE04UuK4iw4atAtBBcaBOQwpJTHGanCfpRCXtLsgrTAo1wELsjgib2MlSXOwcSd2
kobNZcjY/ar65N0Y5P7AVEbPtQK7Jmy4MJPU2DAulz9rZZ0TjDwASeBvKn2fiJJ8
o6JyIl9nCdBWyg0rdmsFw7or5W3KW7E8HXdmIlwN3b9c4qpIih9/A65DnHd8vdSE
9+lHtFJ38hghci3klM/fQKjL4WB+z9Snw6E65Fx06ilelfvMnet0O77Ddu6SuC5c
eylBcWuilIA8R+8d5jLK6Hxe8gM5pAfSkdviTY/QPXw5dCq0Kye6wPJGH3ZjZzaH
yEXzABK+Gkqs/MOWRjA38qgyxrAcTTvRSQjBV/nSc9DggGyeCKbTmAzKhRB2FE0S
+E0vMi9nL9N0V/UkuRxUPcZW76pQAjNMdCx0/LpizdqDICnEJ7C2nFmDhBT1ZWlf
peWV1vYc320eBsO5WDopzW+3qnNXhpUKPOgujceD8i8HYovL4OoTna138bye8Y3Z
nL6xQSuSMx58Gr6SNdN9GBl2WZM6rRO9QawMVdHjAs0mS9jVeTlbFbbf4+Ke/PYc
9TQ3jDDr9Bbb9gxfsdiTxBt6OBp6ttbXyweJpV2yHUPTzMIhRcaxEk6i3XpsjuyE
NX45d/X8VUQk2h7O2RfUEwtKmCC//sp2LP2VmmctusO4VHQ+DWG1UwpKH8195vLk
sOCJ1rIG1EkQCi2Emb3fQmB/j/iIUbLWO0WwjEPV/ZXpKdaxHRC3LFXo1pPlOP3Q
UUiOBEUsHdY0gvI/yqBk5Jc1wrLJddPL1Z8pWqlJ//3Pf7inFniYy2vGbqyku92B
9fK1K+fUy44IQ0QS67E99GZ/ivGmYAqzwQgYZlv47ajcRNrujlA3/mCMDiJXuA4F
9xay/Qnug/nlsqUsNbFkIA829CeS2oy4y7jTjK7Bypz/Ob43KNLGiazs7y6DuRTP
8WEAtWPNDlcoOqUPn4Gm1wAQXTpAVe4+DzH35Vz74KVCQs3utavkOiAdtfAYv0yr
m14JmRp3GQ2+UcX1tzBIuEvmcaguD8BHu2rcINzMXK0mh+rXztQtxTMrr8zXMdmr
aUEcxV062sajD87okksTA5M4DWwZEnSpgACSB6gPCJVo+o7utV/cN7KNiky00yT1
fCNDY8Zy0cHIAgJiqiFN2Yt8H17ufpnVa/byEoH69tPylafenunEKMZ6rhIP6osi
lQiTjvKg4uba0+bgpB6L/yySSHj1t0hyuT67clQv44v5qbk6N1wRn1yZxI9OUGIc
m3+155MJ+nd6zaKO9L0TJ/ZLwtb8x7y4FLUPCB6+GAM2oRua935zbzem2oA+iOAN
Otcq9bCz0qqrz480lot6WXQJw8gRUO9Q/N0ULcXGJJ0u4fIZodcftwEK/dfDmZ5C
8OCGF8sg6wFTRcAOSlZdxwzp1Kp0Gun0DyCTW8y6aiCRXVYGlwJsWUQZTCtcIwfv
Wxvsi3f9Ltb+4JdMr7TGFVj7w6sY2lLye79On/ToyzaDO6TXPtCDPfSBqkOdbkwc
O5l/rZxNJluQZrXhPGjMpgOHAToxTfXQr+CFzCPZ4YlAxPpABgx5DDl1MBIcwZ8J
+rSf7MU8nU70DkpmZx7vmsjpsBjmlMqgwTWgv3qNvRYcwmQo6fvgpNdknoml3905
PL/5c2ootrI9mSnZLvfK5xITCdEICgTAikuyag+oYd+KMWs1hQooc10gr90VfurL
Wo+50v7sD+5RhsVwqX2/dbQ8Cp2pY6X42Hweg2bSetdaa5kS9q+OIwXMsJ/pfElC
JLSFdBjWCGe/tsQUB8r0YCVNejB60VIUUzAoXrvlvsD07/JlaGJd6rhIxFJaqHPR
kERBMCiQQaMtUpVmRVTHAoNZ6HNVNlj/tBIG7hx1GaPAalT0r0LnP7FXYaF6i5W7
XnXt7+iPPE6ai1YJ5qkorgVfd2gS1X3MgXAZFBnfQcHzhiO9DH6dNaCE/QFzcqF7
vE1YlZCOWek2Jy2EetUuyEI54fIKuOGDxOSXeONklMcV/2u9fSSofprwV0p6ohMQ
Skn/1CLmjByzPc0/9M72DoNMfKHsoKp+aFnInWN6uEpG+vedXyk8Wy/GxVUrB/u1
Y1IdXtIoSziRx+G2XDCQrHe0p9kgD9907dFRVmj7fH7DbGPXdwoL0QPaGYyelvzo
hsXAaicilrDT5nb+1Qj0EN/95v6u+BehhNRbweJG9CAenAVT2nnPSBQivD80+rkk
B7s09/SRUBQkCLgqf2/90bAQOZaPiWUl4ikrJ50ypvdJyiDNXRoPVvhqNRLxEIr/
A15258AF37KiyI01cOGYipIcIP8eXLRnxckJLMEh+7qm/0R6Lb1ouoSZJnqUOotM
Q3i8XSNhnWkJtk86I+9zMp3Kw+u65t81yu1BACAd3sUxcnCqQeWStBsfHYbvGhT1
/PUdh736zdlPtikeU5WPh7GvmZsUEajI7mI0eoQXePe1nBDEHs7vG4sEFQJoHDUQ
nf0VVDSkVuEQ1TU7MXyg2RCrisl0ZyJoLy4+O2zgo+Br/HZ19++/U7bLKXj19yL6
B7RK39HeV4lcMqqTXJzEmS4aSFvIy05M+nOtCALIw5lTvBTiUPKXsdeQgwJTp/Pg
o90kXMsKFUY41+5CkBxuzgO6yyc5fF3hVJSSS1aodZ0whELrns3J1008nPadTqm3
5JwLCgtcolOp+B2ZaPYmD27MQDgJuwihVNa5+xOT/m9R4bwz+1x6j6IyLioAn8CU
qQRK55SLxbCKTv5w4+MQxjQVTLwCw1Mgl7p8CnDLBzeeg6jlD7O0zDB2TQbiOIpt
NWOr9XpyVWn1Fb58UUCioYbYJBntLaw4dFoWeTOSefaSICarr3gv8FIhLYNFfsHf
R6KtAVoMhWMqdeMs3BdwvbrXj82gJdWJqS/PoJGj2e9k3GYD0F+ZZZ7TYz+oHi1H
hDaRLFE1cWbXhJpbS5Vd2EIEnZH5iBdsAyXp5+GcR/VB/K/m7ZL1D1VRZ0kYqLjC
6os3odV5DXLy5eTzlulcgJJERmOtphwfH9k3DE52uyZjvKL9sm5Q3I9LgBw6qeOr
e3q50g56AoGj/KWmI4cbco2wI0QkcPvGpN0li8+6EUm07ytDZNpJvFB6H1tDukHM
251/Wpry6RjoKwsXHd2+pr/CkiTY+egDUOVn09UoBVW2h+CChdnm4cNeJy6CGmyw
Nt0bKzku1A3t5kib0tOJ5M9NiAPSzeR3O+2PRUUTDo3lCiQ9cH0/t6/V3A/XEJnZ
vGqKRtxc5KDfPsNRGv/zOjdk9FToQxnc9MXcneTSmBjR5ejt4rXc0gmYxo+RVXJM
XJIN8xW1D1rz4rstQp163QhTG22kcD55Ccs75WMJOufpUaDmtqxwRUBk0iePUCJ1
p5hfoNGVDo8U7HbN5y2dHzWrytoZ70FfOYsoZUfV97YBebnDbXLzoQpLKZVNKdkd
LDbUHh92I3kAC97tQRqemfTcNjiGt4Jx+CqqglcuovgW+hPDjPhc4MFptbnkRdZu
z4hT1+fHTqXr0cH8j5mqXAdgasx/676CHFsPH2jdwBsIrsByj9AhJA+FWSo/Jxwx
MBHkvgKY63iNXp6zWPRs5mJvoUhmjBai13y/rrk4JBKcBOPkFDFoyv+96l1pAtOF
Px2xP5hwSaNtsKqSIJp0qpPe48TEStzrEtAqo2pkElTe3eTieS/DTPdxK5pC6T7g
CcL8xlSSXnMKuSC6qA0LATyOzrONFWOMxtid5L2yqvvJy0QkZYB5Wl+QRqEjXbQy
0krGme7HvuDDLG0OSJSueFxGYyzuiIc9cRoAuXRXR8/2rJRX1zEuT6uOKMJwhjXu
FCgv26vofGPkZJpcCjYpq6TVWWzbH1m1bS2LzRm15rs8sG0UpacoyeQR4+KfXVPL
S+tG2nk9RhUKLt6hSZZ7aBAowtmqu291dkFEG2my8XPLm8RwMVV08Ku3KNEZafMG
znN3TZHkeuck8GUPVX2vlBdh4nHCrn6yAHcvDNGst4QutL4/TsBNdiFnI1icDHVw
XbSKBajOUDaFHpNgiKSKx9ut5WbkE/xDKMNIioAketUv/ux4HjH1H82VrGR8MPKa
6muJ2VkSH3XP/zFm5LZ0vjD5q3Gq6b17sSnk8tMLKOsbDUNMaGRAB2+ggL3+DihU
+JpzfzXrw45dhkXMr+qwMoYW6lhUYm14N4qlZWa1BO1rI/Gbcr9vCigqCvcSZ8bv
/bzTIaWhxUc6tNKenOmQow1PGcMCEWsByhbrstZbHAsYayXRfauS6OMYAwggomvw
rolF30NpFUGi8BCAxcGacDUYe5d5ch4kPIKPBpkg1X8QEQ1K1KrgD1MqRV7PpX4R
h7zw6cCoMbFvhALlNjaiKfySQTIk8P011dMHsGP3OiFhnzC1cS8N0cCrSMKAAH1S
4NehxHHU7STyaIPAL/UY4OaI0rv6xO5LW7gNtjWIKyYvu46Jk8L/vyb9OfQ8zMzT
wFxz8UbuUPXsSVrmaomUTmGOUg5my4wLDuB3E4/dsnIQtH8hFCsqo1XDnOTmFma/
IqrSst5EcgFkEtHerZ3KCy0jg34Sa5HcpvHjc+xlPhoBFpyYnaFWwjGNO9E8w6Aj
Gxq6dj5ZUeWvhKHkExwHbdHWpm91akCiTyJiv3daF1nYN8odbEkIQf6Jd+qzo0Bi
7ZkHOZXeadwrXnyLXkVxwUAoYWN2Y3uNHlIF7FDyKc2W9gUunW8lFdmUMRfeAceT
vY2uD9v5kww2JpmswevfgHd4HhxerTFR/StLpys0nJySp5xs5GpzpIvkdRgyGAfZ
BxnN9NmvklOLp//FOydzSpdSYVDR6eEKGmcl+5vb7gRQtvqhQsRhKq5rDeO+/Vvk
+dPiApPpKvcHgvy1fzoDeNDfgYyuS7Me966gHFXmYJEa0jAQphGiraSjjjWDGzy6
unif2j6Q3PrkN8LfKFvDUgS3NhQE3mk44XPFHor2iu1Bxw2rDofohgXI+FhUhDQb
Hm6NfbMI2S0df6rkUdArnpR/D9xUW3ryAIqlCn9inGvjgWl6BilxEC5KCjW6Z/G+
tlR/5M/XsFE0zr1dYC4e6met88cGRCYe47aHflYxjouXGLVhz3+lEt2Yhf4CoaOY
BOmX2pid4Mnm/cj0B6umzZaPeVEYeqIr8nvU+LOcBOEtBh4oODSbgxirEp4dclVB
TU4uMdvETNWrLZCp0rFcWzDeA59eJf05qwL9FtNLGVSY/lPccrR20S59K3/cCl1v
yTwriDRVrcUAS9IRnxTaA5dX6m5Gk9EqBcf9Kak67tAozMwZavA11sqODy5yHRdU
yr9AOgSSs+qXS560AYS0vR/PLhfuFt7tuFtEzKS7wkYJgjWAIKx62nGzjrPGTAaI
Jh49vO16AC5ys55YYMK0dpjje5IltUTEZiVl/7Qt0LxHtGr1b/xxEIb+iNyv14Mu
ITlw0BLjilw5HL7t3tDtAc1m1Q/J5eT8mJ1cjnCdE57gY/9PiABgRXDjvtMw3V6z
jt+cEGCMmmBCJmNWcLVivvReZs6Kl5+LLeF3e2YWWdFBFQKASSZlXGQmEE2rRskK
o/QyaW+FmMqqnBwpk1UrjoCfz+YIcRk7DD+zcKrKjyGyo1MedmKPc8dOR5viswzb
JAdKgsNW7KBH863ETdHwRPZ+AiS+u5fqabZimbNIrVMrQjHCDmZmRMpK48Pu9H2x
AC91U/BW4CgbNxBFNpMQu5u4OyUW5DPIsyWqcGkeMHOJhqCRoRdQNBebyMnlctnS
PbSP1fvEYlrmaQ+yyrqRyMgXT25Wm1H/dE/nW6sbkOR/+knUcfriJ1xlrKXY+xY8
xehJBf4E1Jc1NJ1evdSFXP6aCWR+8+8Tbk8ZssuZqxhTIVXfSAEOEIkKV0nvjXzN
c/CRuKORm0d/ONhhj2nDddMgYtuiaBA3YmAGmH1ixnXgztltnwDt+VHKKA17Xg9o
WGIGoi4pGzgRoHlN34iaPkStnBJ/4zJ3cR/QVgBInFSTwxdFIM1rpj3D6QKHTQ8g
R8/Qd77qtObVRMGcTrYQCAjzGJiyXs2KKi3nlP0lAo5Ml2QOTnJNUvbpJ9v6DISP
2auIIR2DoBZqJDGNJ0tbbgdqwaZXVoZjf8qsfZ8lp54rnoAl7+KbOp0J6WWuibzZ
X1HLbJvOikj0QIlfxqOWu35zHfq/zwrDkVf+kCpD8AJWQwePZ5R7lmjquBRVtQ3o
SGRYtj8g0yUXiVnTNC0xdRM4+DtF/Ym2ASG+tVrWGU+5HKpDVZ4MJ4Wczsykmd4l
rg94tQBj+JMcZiu+SZ2pkdjYRYhOVZhxKg7Bo2M7VTDInDvktrLkfQZysK7cLcqg
OYqxD8MkgXRrk1OTAwzQmE+dP2wGwOdJwUjGF3JnEuHqYhvkaBrD+imdssufKBEq
aAbPBsQ0nSLnOLk8cefIwUZOhFmNV7iEhwqj9CT1GNQWtMm8GPECdG2ct+jcijpV
9LfK6JMFG90+oDyL0VWhhbZoC2LBRQufUXpC0BPjFfaGMdqAYGYBa4aBeZTsnCa7
4vfThH285RJuGjWb9xGQaZWk8dwhM6PfGy013QSTq087BSdz3IyWNh/Ty4dfetVK
sq6EzoRu4NbcM3f7QHXgrR+hFQsrDa4UC7pmvs3ELHKLokBWfDH+z4MyY6YkTGMh
wkSx1rXEtIvMYYa2/dNjSjY4WY/rXeciv1OXUivwmH4uwbzs/NSvVQaNvwWO3tsQ
YeXmI740h279aZf96DYMzl5uPrgnBqPfJ+UoWvu42AY2Ds6xH1Z246KAFumOh+xe
0aJhM5a0HWpDGEcRZDxJs641TA74lDz/DWoS+K6JzbEnxL3yRAoZVvaFco+vDH3g
iWoWZAM0LCzfmPBvTTE8q3qtr3/wyE/sZn3RoEqfgv/e3FWiC1VhZsyII/9nTYrJ
IC+PJj74DF8ag0GDW3G1MfnM5YIhbpSA5hLcNh98b4wv8DqxRArfLtCIen25/oBF
WEA8L5cMt5lzgUqKdlqjaXl9CIa2bHTyKoVcyg58J7ZcbCxFrO+ipZkAJftRkTZ/
pXaK+VeJLs0UPWX/UTqeNCQnP3Cl5ROY5JNiNYJtvbssnUo4AFPIQcTrhL9Ty9xA
4dup6KuFIEItXHxErLWaZYWt2/PrJwNzkQVSWwcKfqENiU2Vr1Qkj7tUw/o4f44s
BN5a7OA6800qzjye7fRabsSjq2A3TZdkhe21lteYH2RwNdFODFGbLTqSkG4mZI6s
5wjVw5DaVnzUU6qIzioCwBJ1nIrFBxq2RTjLDPlxx7QO+dQtUqNxsMK2+KishHkq
aBgfz2CmDE1d9WzF5l+Zz3GlfjYCzZ32JuZFj4fyJmYzeBapGDS6BHbMW09PVK7q
MRv/pbNvTq8Ausx0M/FLgioys15ai67qRf5QALV35WR3vJEKezuujfA0hjFl93Nd
vUX6ctS8zlWCQ2kOxN2gQMZrecE/zov/olBnct4eoqYLM02M//uhh0kLcQeTS25h
bFKXedBPvgIeS/YYrFPRbRJWmuZgC3pagXmgxefabvKSeWUH1pdGBOjeTYpoYVYk
UFhmmEqE8WM1gBxEDwBDjEHu2RjDbU5GUB1xseYgzudU9mKnxLLAIzEoYueeo4xR
3iQn7tIwkNQf9CjW4GwCnVaCv3ZYvqLX1t9F2NDSlcqCF9sb2o8ZOQPo3rSbqzYC
YSAJJipiisWeJk/hiHim1CZJbgs94ufAbEl8GT+BRT9rRrjuW1vX5cNzn5LgulPE
5HO7zw86qYPPP/tcpo47FSlgjsNhjK59cGRAVDmygFx5YpjGWlSWqTnXMBcNiNIX
Ws2ZBRmaQcktvB6FVe+XHCwNvT6BdjUqU02RvbZ6akc6z3sc7nB1ka0cz6h8fcv9
VTGWouzz0Pm291DXCO1jpWtIfYBHjABBpk72m8ckfNn2PPY2LmnRidFCZQEFd/YQ
YMrL1DrvRGdZwqQulkbxD2qQB1M811QxJIZJ6Soz68akmOLbgfiU96wtj0XD5Day
ylEprEHICxZjBeUpFwAaAzFPET+lvuUYcJAdVgEWLQZuJaVKF83tZf3BxhsAFjET
lV/Mv6q8/PVyutZ9Y95pyIqLvxgGadBavjZ6NIBWxBQSVH97Vlt/PIdb1AirQNMA
2mPKOIms0mxnfSVRpWIHN6JlFmvITMYNfz7IUSMtIRSj8ck9q+HCoQPaDkO/4Hl/
jywB8UiPAb6w3osalPqoogbHjoduBNUYxu/hNAjVEpt4zqLoXsnkmk4mhyMxovRc
1tI/wFP0qwyw4/gl4j4+9oFBWxb9TpgPqG+Ty2kD8CyUHgeoHcwg405W/ubiM3qS
fXRlc8Pjdzf3Fbz34LvHaZ0BkhsnDvGQMvMZO23vizEqr4QAX7SRFB08bwhrgPcD
AQt23fINCVg2F4rTmpuH/XmMPy08GXmjzLyshqadCPle4hetQ0vSFNpAGhro+Xv0
OFFmEAYXmqVUtCj0f4M52kXDWX7UJ3cL1ouLBrwqpdyxGHplwfhOMfjxwTh03kb1
27JHjGl9n+LnXO6fJfRt+QzZDacWWlEJ4ymi9PfGK969CFCXVV+S0HflXlMqxdBi
n2eGS5qT1Llwd5h161aPUx/8fQvkHR42ISgGBB3cp2o5RFVtTGCScV1YltdzSgxU
jcu/nls7VtD8O9mbxvwaQIzNcRA0wdxKAwwPo/xDdqWkjZ+ayoBhpm1cCLdhIkh/
FCnMvwG0uhB+knGyrwambPocH70PigygCzqzy3ywNwgv7jmJ7FjkflB1Aer/gSEe
I4vwE0S1/ttFMi5RjxYz9H+7U7PJK673no8fCz6++ZPFZb4oG3t9WFGUdESKnHXk
KFz8mfC4Jkqd0jjBEGcdu7NrxnPoEcza3BAdsIpcbq5IEyJkba9sGxw+YIJVUSKh
JqSWCgor4w+7Wt4G/8jrNdsUmSdf7gCBgDVdVFVM3rUcHu+5YlpYMNxjhhpiEybj
XluZo4Uzyke8Y8OeGWpJ3rqphVDKHO7wuUygnxiHLLqU+M62iVot1/4yA7VIOHAf
YrQ1VAMt7InIKFE5qGT63bYqzWeG3EhqPfZxWebPUK7Y/4eW1uxZNyP3hH1zL7Q0
0qGaBOo9UOSG9vmzYNkcosDTuFpNJzoKjCC7RS9PnRq823LQTQjFO2fuBzn2uv/z
ShMWz79k6vFCbc9f97fhvm9RoRF84A9TKZiVs25KzboHMvR3tfmTxEFLAoiuuNEh
IwP2G2+jGvklxbu3i7ta89sihUNB6qULRhn+CxF8vleCGrIPHk9pvJs1Nqy8hGrR
Ro1FjPI9E68+stQP65fnQSPEQ/DuWrxe/Z9bXVEfqlb+xBzuACbChz+0Wd+vvTfI
4WGftySBY+T4u82U1HM74FTirkQr7vNugCcIhqOLaQuXnS/pjRiUiTSKBRzSuEZ4
BLvllmS+BgaxoGSZoftg1L/vLKlJ+ANj/3kue48C+1cMbMTv4aAcl4rTLk/RtnNT
vyzpBJ3ROUYzZKQTEgESmNA+Oc9EIT1dsGtYgFwPEfpW3gk6eujVyD4l8pKE1958
OQYAJBPwMMcgVvPgpvB0OwRVSkuQ5e5XQKv54pfxFZDdo1CsA6ycWZ6wz1cEsm6r
7alee9+RvlXyq/9jyPSNHYWDJtE/R7kgMA+ZJS/b5B9wJUBHut15HT52Q2rSue9b
CzjtQodB/P/C++YCDb2tFMMDfygei4Or0hsiE/F8vhlQLuWfmxjDKWoIbzR92Kbz
YiulQMfhUt3GC3mR0mDQfn9x8wdFUN/cykHJLwdhkdhPCSKBkx+vYPOmlkcM3DTZ
+Yc7tjFgud4An5B/2U0gHNXZzsyAsGkMIkeJs43QKiXLWamoG+/8gb6bWob3y3e0
Wqcd1gZIol/tYu6cOvxE/QF3HQsEXU/fPMFwjEwz/J7maKHdYuhhRFBsobu/GWd6
U8LPhAspQfLaC9RjWFikhm2b8HsVHJI4IFECyb4JPpEUOrw2m38nuEMBBjXkDSty
BAoETS4dFnuOwzWo4RWAHqGSYMnVXgrnqFHJZrYWX8aawnN2QjgfphvjKJO+/EKo
n6DlCIMgdCDlwDcOfw8eO9TS/I/fu1JsH651zyibWYxlH8lxw0Foq23kGjhAjIn7
YX0zEscdDOOQ/V80L5hh8CTEI8lIHWcJj2g3R0p9Pv+vIHMW9fr/4GjvejhTCzbf
egE3osM6MxUoKLl0VO82EWnrZc0JR8ZbtVUHgPuOeS5aewDGLJ+On0OGh6dBUdxb
7OGMLBiXdT25+HImfkS2wlpLFY7J+fSFrEYGZAKqrNABhMC5BKoBJeP9dPwvBE6v
hhpYKaE3mkWlIGck82ECDm7P5t0zCYqisDpeC23z/eIkFmC6O/aX2v4mbakcBQCW
f5QsviX6i00G5OBH+IexYqDOoeaBfb/fhQ29a+bPTLmwVUr39GfpmizjWEueAXDY
WU+64Y3mCxuyFFGEHFzRWX3IPUpFqrKmM+7AnXsWRLjs4N5WEbeLxZ8w5X4tmkCC
BCu9ttBmJ8Z41hT9FVSCkvRH/Z6IgBMQIooYjtYzOoIkfo/GCf2Zv86aXi+xvnkz
Ap23OofUVRDwB1NcfDbWiQ/zhESV7U34Tnv7ApDaYxPeZAEomtGBPlQEajvnOYae
oxZmXhbVgb7K3weMUFWma5lrUGRAlDhkf57+uuvSTqkg9qE8tYf6l2T1vy6bk+jh
3ahsBdYyd7sSj8rfnKKSEUYvmYqmnqATmSkGBHPdh8X/VIcACJ2J0ErOqkZTrM3C
3PQ4VBc8YBHI7HPxwfmCkywBkpijvwu1or7Keb1zGw0MNZ9Et2kGXWqoQOgxlO6f
A+3ytLYsZ9dqNQOuCwbJDFWJB7LAU1L7AQT6p+8iWAIwSU1geh0mF1YOPcyeOtmf
pzcD61XODrPZTfzRE3hAslh8UmcdOaSn/bP3vN7zCbaWJvLTDCs1HTyUqbyUZ6ge
KqcCo1FvYxYXH2ld9jJ9l2+7iwmqVTfji+AaqqgTlMITtwb3YlbjXIlB8t9AE4HM
h5qFV5/GcsmsMaXniHFSwIJtokbuTAIGlCWRX+Zt0fZjKO5eO/DAzB8LmytWPpbA
HX/zvzEhnDg+5KVMMxGB7QzkLaHkkacNMMPxcSV27gj+goMZqWJmBci2eUODGyRQ
fUu66hK6J+8dyEf4Z4keFltdfw4xrhW3hwiGmqKhHRhizexDJQO49H8vzzNQawit
Ftulwk4tNVGuxiyWLSwjMH+vT8Dtj6zs99Zsq6FZRa3hG9Z1z7i9vMlPdHBxCgHu
bR4Ee1EwPRO2V5Wh6nVmtqRoGoI1QdyieX02z/2+w5C0OMuJ9ooG8DM/iozs+yTa
CubZvPUu5CiVqKQpFaF76RNR4QMKFv0V3LzAnDdprBQFIMIGqkNamDhBCjiH5lIV
E9KtlHRCpkIzFOWruhE5tS62FRqTlFb6H5xkVKkt0Cx1wTfmqPe84MvRLnIlMMdJ
3ByYQlr6ww5jNpiOyZQI64qiCubdBjq2ab8lXp7nLb7tnKh9tOK5yR6UQGO3MNBv
vuud2fVC9+2b+WvzGReLrGnrU2zYcRK6cexozPrPiHHtueg4pw4SPhHWUm8EoLN+
jyn5BKIkkblvz22dwLIIHoTTPEHICI0aaIoEVUY1YxYiaAataT4G9hUilSbvG7ua
P8cr28wFVLqPdyIuY3w/tL/yH/59KBL3yGNGbLWwsbJRiydkm+rMIrDjLMKjOx2+
q1xi8veX1kxRlMv6gk9wp+XRKZCYSCaJI6N3nwB6wLto2lIMSe8VH83E3V8/r88u
fiE7kHVqX+yn/NaKEcOT/splKHkWlOqPH07BqTyDKxv7Ub/Pv8bzK7zb6+JofWb5
ZMhlWlHHHF22mh4f4TotW8ZZJY5Ilmd2aYs5reTNaHMAVVj8ekbdFr8my0MhfKEd
T0+zl7vwBVFYP0beeCPtidMh6xznS7BxeWZpzRYJgB8LF1UwyNtzSrmuvUxUF0G7
MkeUTsOnc+W3R77ioMl1hFFLpbugbcI2cvtf7AqFu5B8VA4FknDncCMFHI+ptI0c
LT92ah1f23ygsb1EL/ei0RisZjVZWFeTGQQRNORophSuQ5AQYOnyQSy9SrQzrkoQ
XX5RM7mhzv7IZsqTGEWgiioQF5FZ1Ndn5ynWbekB3q2u1R2VlxQZEZXPK9ZO90Xx
/+STxvpgr0kuShZ7Wk4H+NvYAGqHphXlPllQhrcUyvkKIlinfNXhsNRSPWAZ52uY
hUn25wjRZuwVJ2iAaU9hepBmmfhHOBdqd9vZXkhTvgFlCERq6r/Kb6dJP6HvIftB
lI4Y58ptpHVpxNdzCDp4gKjwJh781wTtJ5wnNWWH8CEyPWqdFPZRs+Huji61PGT3
5Df0c48hJEn8R5Z9qM7fHO0SG/Xfess3VuCVX6t787o5tG//zvFi4diLya6+Ad/6
nTvGNeQ8MvzpGXVQysWeuAa6jad8qrDlb+h1sBb13JzNaPGiDb5zHQUzqkrsCvM1
qM1MY/nkC3sdXUJN/G4X1TpNIWUzUUlQw7rVxIxN1M18y/pNgBwEGFPFlBf1mJ3s
CaUPBF6akg82/40lfxwPTFTfcOHc+TwAWI+ZSJM5BTzMspm+FXZ9gnhTYHHebaN/
vlOYIxjifY7Vel4ON8GvKIPyVLv8R+FDX/Ob7r75w4EwDn8IzPi6SETV/Ycp1nkp
sXAka4m4f9h+W7x0Mi0q1hRWPg5HnsS36gJddJEDG9j8lqP/LiSzSirrjcjc5H66
Oa/YpAzviP6Q6RUZk++lvWxa7hDBbjizVHgITcS3OtslM0EZLwTRpI7hVT7eNSuE
DbS/PmEIdmn8Rp9/OHd9DAvA6jrQ3N6CeGStFgWhAlXfAJg9vVZmEwSbQcUF8y8z
0B3Tu6HxrgYRLnVamaRttefMe5Lm2AoPEvxx07s+FZJ9akwALG0iUPqA7SYnReHY
yVa9kzZfsLmTfK/0E7Zf1WzdgC7UF6QK/NLp0vToCKyQITxgSCLn2COZVSpaTzTa
+5TxuH7R0vxHvFhlQyeCgXU/uVhovji3tbc4165PRov0n9yOQs1BoZTPuWHAQ5Bt
JaPHTX4kiRrTVofF1Qvr8m+0UfH73kVR1OdW5Ar2yykzkRWqZPRs3ZMkoqnzzvKk
0A5F9Xy2ifP/MNQHgw40kb7n2etiMrVlVaixmoqF63xTaRV8z2nDPFhuaiQS/m1Q
KYtNzhqUlVYcspzrb3YH38ziKI3/7lupAnQQdGYG/6u2Oq/PDvnKu5laiOt2Y3bk
/TsQ5+1LdeaQlbjC5RrcfBqn2ZQXKUoyIrISqZKqXnLS+FxOUTa8E184NH2BTsCz
jN+ldFC8wndiNgfUdHq5Vl778hin+Fw59aPUxpY3N/hSpnbflhraXqychvTZymXL
rzVUQXTZfj4NKzFbySWnRrsgyFtqYAYFAFTdO1vDwDm1UFE0+rtftHUxvBXVWMyB
UbNMEWUaDVI47qns0tnmJFVQPA2gTjpjz6yCqjNVSJvxpu8BMQVadfVrnXdUHnEj
3kXPoDJSnONimBME1u78BTMGX9tbP8eQ9yHI0nqP9P8at2X7he874n1SUaSp4mUz
OPorJe7ko+NuCoUEHQHjQBOqdYHLZiITCfVIDky7o6JL7xMrn6q6FtrgEsgcOrYb
vTI4VEeilD7O1jqGzZ7WS3xYnObcJ9+ifR1ncIS6t8BoKT6v8HGafAcXIohdit+Y
hT904Hz8egJBFoY2TOqRSlgdTuFFa9sAAPhhxJZDS5k+FGuMngrub6s+lBUdwu5E
ckySzv42r23cxSDPkVjqRyArN0VRnuoe/pMcUGC08mNp1I4rsveNZDU+Su0eq4MD
hjHwRyyb5PI9mhG7KG4azcxu8mF7SGnvTd8mSeyBrEcEpS9Ztv9B90tcUPKDN2yz
oUXSKymNV1ZEiWYoqgw/vD80slq+OG0jF7MO4q5+0nyHQEwqhVtQL4eQQrg2nUBD
DD11UNkmubfkDvbElFkYw/h6P+YfXn0iat2FmYpjS0lF7oKosxSXKOjLiP3DHxUB
20994cemYqCDZHSZWtHZkPMvBiQuvwD5DvJKDn8K83mOuOT+Zg5ETAItRMzLms+4
q5GMtH7a3veD96T1SeoLbE34U2ZuWozqGzwt221GMOTrVpQHw1uthmMljzG6K0rz
pEm/cMUtL/QpGrog19AVMH+GY/4ess7tr22ZkIZFbKNrdl1sBdYQzWAYHXmWy1bq
YaDPTmkwCI2qqwZABnhGV3OSVAbPzNAyfV6/nk1J7IiM3jsyjnk6CO4tgXmxfJMJ
zsDop3T+kMNkkp7/YODu/l1/YK7NyJsMwc1RtviKUhriTnBGMnuyrU0p0Y021oat
Dg4uegBvS/FxmtB1Aw9T/8C4ZLLV98eTR3+r/BjGIwu31NoAGfx+A0QbP04bh9pG
M22NCStJnMIHeKwpAp3v/ws1lWjv0NQayPu+AsulXcgXtBYEFOGWOeUP7mymxoen
gJ6Mf9g4brQTieLthfKNPcgLM90gMfr42E9hpoNzPGZBUrtM8MoUNbJ+fIBJqgba
OSvB+iiebrruZQMNKyRE2hGFKmz7b/0O+Nz/VrPpKYvc0po2ACXxzLlWwrlLJb/G
IFh2Or3lLbnkMl1cofPCJek7pIUCJudEOTlwv89Gozv8ZkUcLTQ3U9dxR+XNdyLO
oInKNZ9FvFV4S+X4/Z+UdHdyML4Jn9OyRg1ljTU1cqOErlkI2LdvQSyumsSznoJV
fYLbq4MvOs5VN6S4yVMLUxJrXlUKj2o622tbMQfAClu5RotBtMZ8jOr5e3kby3pH
5biyD4esDBU8CnSjEzubLKC3palNaiipxjp59HK3dnbY4ZOXAmX5I8FqtE00JRhd
p/A3Ln+avIQpx7cQT/eqfcrjHYaqUl2/DYPYOa7aUOJ+6aHYvFj6/NGC1y7CyZzp
9OaFYwe+8EQwYjvsjFiD7VSiaWVMgWzFBC8oVTWfrDfdee+Ro9Zo/WuduapHRPBx
Psa/ZkrNzv00m2bHNjbkXPQDGPfa1XqwYUISTWLGWKQMosWsmjXnOZK0fnl243uV
hy+de/Gqq0aIgIF3fiqhZnXeuo5zNH4akq3hvZKXPRbNwLdcCtRV6e8k4HoVwDKS
H/gE4QIbNLNezh2WNGSAS47FQiTihSEINU8YaiQWo2wdE2qf8pRNi14WwvNSO/8C
LMnJ7bRZp2JubsN9WY7DQja4IGmaUSK+pbKdi1zq+vFcDUeKcey+4pAhy+Z3Rfkj
ymfr+BZ2F6PXXD/eiejavFlhcHnE+Qgz4McA2HLI3Ez6mjLsqcDdL96ixnZNogm3
pBfQixX89TegPZRTxufsKPcHiSJ1pIuMqnG0YUQLs00dnpLeKCL8mWG+1hTwX208
rlXD8z8LgxRy/D4QUlCcbnet2k0pslg5ly+8dsYdjPRqTK8CGs0QucrWWPafUxfN
gcOVyDavH5ElSlM7w/0xpFCs1g1WZrOURXyFqe2oX/3A+J3wDNCxH1QNA6Po0KHC
v87yNhDvYk9eqQ8kWHNUa6Cq914aPcRZe2NqKwBxsBtc4DpDKzClNsnt43WvnKoA
Ern8aiHU1fFB31BQmEAnnnt+SXB4wEzVIqPP3XcpPPDv4hxgkz97Gn1sjepf/E6V
OTsrRQH0ILskPDdu/s6zr4ktqS7usVH0jIQoKaxw2R4fFBmKtNbzF8cNBzLpVUuq
CJlqGG+U9gk6i30FCuf4p2N1jt3RcsFP4rxGUFsQPluHEdi9dIL8U+QjT9XUDRf5
C2JlB/MIDbLTEydlVJCylTixgz9B07OClVQ8GWVDwj2crYjPz+l5h14HtbixhvhL
6cE2aQIHhplWRdPozDEvavoHGd5t8O76xR2So5LoQrLtA4nq84uMMZyYza6WtKZ6
EdB/GpVSQSFJbb4okO+E4XvKg2Ml+7/LcLuYcS9jc2sGbUfb/DtbtPGAMsyr9W5i
3iqTa3OiG1beTcEAhxwy9Zac7Ta47wHfbvTOrC0iYcecX5JhPe+iea+QtesOYRUB
vi5ESjrUDs2VN1A333z52SH2IazUmcDbmvN87XtgmrflAEecCs3fFWoFm75+Gpun
HAzRzHrO5SNVUwIR24LTfSAcvUZg0A8dW7xnZAIyheQgZKejNhpJ2X626gf18EPL
EtB5qWdM2wz8FWJudIuC6YlxEhAkf0ymBfg6Ml16F6GJD3Da8Yh6+ik+47NuW9J3
PIYr1tqx1fWt5zCJqNrMGZQiSIkHlRVDVf9Jxp7s1Ips2KOc1sl5LCPVYz7KjVwD
2sYKIqdpxtdemkazc9E+5ESBH0O+GZ2MBYP0ritjf/YVK2X4wM4amSErZo/IML+0
FKCWK9JE1+OD6ucKrO9wlHEtRCRGZlGYabDJ+se3UtXOEOK3jpNby1/J4BUzHieL
Bw6HVwwkCVw4+iOF64Jx+CMKaIgxFDxAc8bpnQ/jyQkICCbmM/v0aAP3SPJji671
w/5tun9gDKilQGcA5+OVzgWY37QsSVpy99fx/S498fXwIHesp3FMCw9mIzJNGnTs
Rmf5oQqjk65YaA6uKaFDImiB0tHv2KvGuU8orrRI/EzFGI2SKR8ICXDFDkr8aQrN
m4IqwHooSw6nrpUVFJDOsTsetwmzJLBkVw6QT7RkSbR5POhYL73DO/Zk0Y38+2aD
3yUdmu0r4DXcL0mcjPTeuI01v3xyKwA5lXaBNjAUceQLeoOtoJXtE91JwNvU6+hA
vhfQA+fenWmwhKXR6ExNu33fZETkU5dOIzigQQH3qv+nJ5HXYQinCNtFHAxZSF+z
nF0A/SrN960pyBOOC+TcNNVRcslNMh8Gm132nxfgbhG01Ogihsqy/f93SggVSwnN
IiCYxWR4HdCtUU9/EcMs9FBmQr4ZW787Qci070IKXfEh/Izfc+RzBbx3nreB0619
1yppgRiKVsMOlJwiVKjCjjLQPTUl3TQakkxy++QI/I0lY4xnLOnsOAgGhTyVaRG7
sBaqndLatIKyX7AncOLEFgQyfVp9WdY/sY7haZIB8o9JA3dqoJYW/f2dryo59GRZ
KYAMKJBkepnmJpsyUHHGzg/atiLs0rw1WkyRIVCLE2RYC74QnTFYJUGmUA0KQorl
JXoKyjAomxciP3o8u13nQteVRc9igZnm3S3rbCZBvvUpcwA/eTZCfJ7F4xPUDRAo
4AwWekQh/EnG55uSk6aSlEwpEq86DixDFWUOccW68LWLYcojjCZY8oFK9E/VXVR4
kUpWQcxhKYRASlsAzdUdpGVPpCozEd5YOa+LfBddUdxRY4Xv6GremczGf5uMIQ7+
b0ctrQWMur/nkdF8AggdGcl9KkC05NdECkKaj6WlT7f9rENhd+Yr33uIetb7M1sG
5KsQw5BiomvKTLILzwT3SCk2Jwn3OA9wF5rV6FI02lbh53y5YiybB6rJXt4zov9+
cx0qPEj2sbwhQLngROZ2XIPDTg5siktzjAWJcDpQBl6wrmhbfEZjLF1ALKIGB//L
JFFud4cTOiNn801FlCi98MSSUn0pBtAlSqeRp1jR/UBuvXNaAD6GY47lOl7yf9Ja
6H0O6vv1h+YWG8rzNrkEVrxGHImsMQU8NOlezRv28vC20X9NI2bPzZ8Vqc1PL/PN
oy+ffdQCZ/xQXV49kgo9f34LTGkWzuyVUTHV8utgLTaQ6Ji7kUF4pei3jZEyKOee
wWqTAe4L8zQm5EZl+HqKbYgpcsdq3c0di8u1p7P37cu9CvPPVAim6KPHlnF8FwVJ
P+OkGE4nPOMW7tXSsg6JILaqbE8YnXx0YDVGST8DQEIcox6BYyRkvGOvWwmYXnxE
i8GCnUwk2wgSOpmicPITy6sswMhQN78L6k73qGjiRetRUc5X7OXEPVHWQTM6vjcC
K2/cOop3T3wv4Nz5BBJuRkiBntwDzPPj+p410ZSk2VhtebHiatv0wRGyjk8db5lM
EoApnc1EiBM6qZK02Uo70POQ56tEo9NwBS4j4UHe7AMBfWoYHWjIGwEPbPKpsQWA
DM0vZr2SlFcdF/17Id1BG215HHpoSRn4mjZBMO6HJNgXkkOfUyqDpnc4ay8qjFle
O8E5ZWOOI6nUHmEejAMyZlyOPKfCdxFfj/6c+rbzmfeWN9ZTbzuivMTliVle0FFb
rG77BUrY1f8cm6QS8EfXyF8vcrypMKO3V5TvyY7vBeubuvOwKrCQR+1lEul+6vU4
7wHJ2WKXxhD//Z37EKJ/SXSjtBvs/JR+Hsr7ObNYXRSmV189GSBdQnFSHcC07xw+
e89RMli6IUV64OJh9uCpB4QjHLgbCoEb5IHkjtf9YY2yS6X+/PaY7szXGE+4JgWN
LtClf4eAVP8wUQFtySS4XwFZHARJKv52pyhGx4CGxgDAolafPg5or2pmN7G/FTpj
D+EbJOsJUN4cpYmlswvdFdkJqrfwxUyTd1eeuvLDi3s0tu51fnI/WKJ+P1f+FUub
UlYsE/1Cwr9yf+Thh73+5wPyaYSX6EP+wnzCVRMc8asjFRbReUj5c1zoB7WAz+nm
vWUozb71roOyhxAEwzVBvNvC0YjUNoL61jtr5AwWK54qTN0Efqw3+zHClfND+0gR
ynAQxMWD3rOFYsl4EDr+LptrFsmQVynpoEWOfx9H4KAiW4gKX9Z7Y0ypTSSt1nTr
gfUdVKTygKOE0o4xtUPrIA1G+1qMYG+1/TvTK7sAO+59gX10BoMwYRG3bpJDRUC2
ZQhTqcaJWAef3xd68FuO4bocBGhID6FN+Wrnp2fYqntdT/bIn6OYpBj0rP3VyBWc
R2smw1GsTHYFA1Rrqs9d04CkfGFGHwDXTN3y39S12fyzH9SnPJQt2C/mA8IlzE5C
M+DAy4EZYHUNqMVtZj7gJYJ2iZ/MzjHGJpQflOwbo/OM7yrAjNnyqIZ00YnI9lCK
bWosj15fICsJLGdaUvKRIXMiYbYBsqsOiqMdOUXO6E6BLL3Jcls1D8KEcETPIAM5
kwYGtBvkWppUy2bGSKOu5yZ7XKrSdNvqtaZRQYYb5zojZ00f3jGmHPumB3KVLf94
b9/CygmkxiRkngXLi+zCYdW6R5QQrrTUM+H17hKyf70bjXfI3Ex4K8xnFjkZmbp2
2AVRgcO69n6a7wifqTGLgzzjD11c6xLtj4sv2P2i//uMZOpAwOsHtEuhlfcYowG1
fhpHBhZUq6wynnL3OyZQyqhqyvotTiLodwH1FGxLylbuvXABOhBJj8nFBI/+pn6F
GxiEsk1jwUD6TburnPI4y1miBU7s9BrW+/V43rLKoLB1dPMl/rUW4hXCR7VXr3tF
mseeIZ4kPi8nvt+M3nhVfnTqUl7B/ShJyQk/YL9BjmA0TR3Ppmn+Kmo44xQfm3iS
vL4QFq5twqWhSe9w5UH07jN/5c15lj2Wr0IZDd5doMKPUqb5PqOsCY3ZyB6j2WPU
0MfmCc7MmwRrIsraA6RG/+qWUFg+u1AWuOlYpeDHugq9N3UIfLHnrvElVKdlPN8w
NNu4IW57e+Ner7JvQmdUSKCZw35cS9C1/W6UK/LQL97yyOzkYrGgW7D+Zc81ktJy
w2h/b2iAOdUjpHXQRxQQ64P8ZB3PruOdthzNLvJmDSq/aVasPEzluYoRkkb3+K6B
0g4rz1b78WhycPJPzJvyXFtMX2QWBgmN7qub9yBCJEQIbcWZrOHqnuJzyObaSuoB
u7mZDEi/OXK6FrIgvKIXvlZjDCrdYpTSjPbaiTB/NCvPGXEVATK3F7z1EzmYpgnK
c+Ge6sTu/NzTosvh7PHRI+xEwzHavHAtkYiIA1Ax3jED73HO3NBTwNNQWqZX6GKN
WCqXhWjVIFR5p47MaJMji/WaYk85h61qIXZhprFTA3rIlHK8N3+WX8h+aSyFfmQC
/NV4xndEcTWCRuaIiC/lq/s2D+TE1VtaqUehYf1lo5IdIcfwRYurhpTs6CUE2NgV
o8hsXgPPHfDpxQag1ZwAu22EIUjVoExqr6Z5T7lVarvOLr/B3XtrHy3LOxUU2Epr
l10pMttoLYBJ7nmVsMZP+wYAp4NwM+3pB4fdSPCE1J1YpReV+E0mO4cU/QGlx5jo
piG9AG2mzbN7zztKl2g6zC+DqJIyRjXPwROpeU7dp1pkVHxG8ueiBu8/exF3P0oH
m+8PGLAkRCQf+J3K0O8Qy/y+hy71Ts1+wHoPH+joBQF1eRth0auYNJBCSML6euuL
3J643KEYYlAigN2FI/P+2a7PfEkluyZ8ijYkJfoXnZ9f53Jth/tatKgdh6EmOr1r
xdLzrFIZ8bS8JDUYrzGzekGsCKCbaLvkUy3PFl/PS1cIG9oNHvns6soNdrFnhmhG
45n6Usqw63md3Y/awhRSAvb6wx8hm4ML6KNbVWgPdoa7MufiHT0cmJp8I0tSJ8Yb
17CK8aNOG9ULH2qWxyNfK8iEe0y6KKwB0YxhhdckblMWjJ7Eb9ZdYrjv2ixObcAZ
Y3jueJZ60oCu5s9iF6jNFGN2hFLpWuNQfIlpY4ZWbQC/CCwEQhaBuNwNgrar9kj0
PrjuyWJuYA6CWfw+NWRUL/3VNonSHGTnDaoUbQ1Hi+IdE3JGtcxzWXPOqLWiyQab
K02cMlV8UST7wMg24p+ZbLAGjT44utd1iSv9AEwxIUEfn8vePAMmexEsDPEr5jv/
1HrvLkoUrZJUkWxvUw8byDc8pA0z5AXRvIfKbPky6fhrSBn1WGhPFHuPDGkdrSaF
Cos5NL7eekFPVQ7GuWoiqR8JhD+SosPt0Llq8YxjXo0msSRkPRW5QtHG4BEyYSQX
MxjiMMymWuDEXsORjAWSCfAOI4ko5Okfq2Vj35GYLEaIgs8CjBKpWOyT7UMQLQWe
UU5jdbsBBlm9bjAY4OKQZtGWtsSVgiXIYpqFO0jl24DmmJOafO1/r3K4Dr6OgNpe
6XdOzXksG8SWyPkQmASb2uJnQUzq+FJcvK0PStpHkXIrC8GrDHnYOWzkGwJwHnAQ
V6IiymHxDQW81sDzKGsD/tw35tqnk92hhNZHBDiCGGT2U22zkBSekbRAi/1WZwtd
LHn/89ArYa3ZNYzrGOBRlVspM5vsOKSVyTZFtLh1BYnAb8O1WHE+UQFs+urj4xBO
R3cGXEauMJM7+O1hyMmKxac3L4QrHr3E54uR3kySZOePdLiH+tkuBxxKsKs6uhSH
stIZVOMxRga7lx36zBxnHJs63W2Xht0Hi3rQ/CQNaev9bDNntM++jUb9ylQE7M8d
9PBgLshQuyNXgZrc5IXRDLibFs4tiSaBXpyZqW4L2Dcxev6gSNfFafU/eDPW8frx
zKWpmf7PTEe1/vIP5wxwkq9d1ERz2YxSbr2UG9j4aBkuKA7ps40OrkVznFNRBiDa
LS40Mq9p8WLr3fPyEIs+X1MOq6X9lb6uwWOrUt4/RX0uxS3CIxu7cOZUqnRioxiP
qjSD5JJnEKfj9cM0Mvr7eHIylBfoz32gRHCn8PQ4Q/i77h+iW6oaDMlKfAaCMtOV
M70R6yqzfyqhRSooDl1L/rkWArJlK6ALWFu9lmwFhkZkwiKv0DO9nbRj4wrZ4KNd
YGAotiu+ltP969kIMxY/tzRUB6qg7D0s/haSzb4wqsGvMr4Xi9RPG8W6aQWakPfT
clrSBDoIGg1xhLHH8qQ1YIiW3yQrjzhEmE6foIznant1cUDv1HhNzDO5zT0M6zi+
O2fx6ID+LhWEOXPA66V0xHlL2LJYOC6Dw6toQQ2NU57pc23DDpP/steppY6x58TD
DwZMhlIkRrPMTcyK9eCX7VbUadQ88+Za/c95WSTiRS0kCOkm/l4xwaxsv35pcGHd
otnIa7Q9C0RL3ieTMSogU0PMOqfCPZ9Bn0fchylr6gBzt19cfuDT+WgyuMGQ1o4Q
fnzYKuwUicMj1Pjt3Tuz4NYUckdNhu8ohs3iUOP97OLtgRdvWII289JgGFcedwL9
HJkLbVEaS37VKNhLUDkW9pw7x4yxtpYVQ6yM9S3rCSCptCKumQz1i8So9AqNc0RJ
xbVtHT75NntZosZ4UrH4FHDqr0/+t6fSa/0PMfD6/fxMw8PF1Hc0QdiTjgKln9nd
REVFXMBfELinU2Qu/CEaamYklPC9hUB9AFfpXJsbqB/qKYdvID9cLnT28RXGJM/t
IwUgNeJEtPtrXstgUYFxnvy6i31B4uxLzjpL+Pv9F8/KT98EE3hBH6AvPlbnWnd/
LvJPd0UXbYsvKwHG0HZRvTH2D64nWaOpzMKd5mVjgp1bKapLQN8Dr+a74z0vyv+w
Vai5Ann/p7GKlWRh1Q2W9DbKFLPog7nPmPUQSQiY/g6LFyycS5jPtZBFjLZ9uG9h
2DRrFgVr2aCGXROWtHzU2D0niHcgBOnl1rmbjcxz0S9LAfFmVZ+UpfMPIqK4Wfm5
dF6zmA0qiyI4wClcWKCFMUE5VFwnjp2u9V8jw886cRjw+ds6CXwptnBUMQSGTZWN
/6t357EU5cLSbdyQBjCNfGrtj042oBdTGow5uoMYzbA3Bg0RvxpzAbumddqCIszD
KF/vbLMUgw+LIk+S8f/WEE6aEN00NhvwmpA0W7DMUxwJZskVpLPQUCkpq878sSPU
KPqqdD3fBh6NyN1q82WwgAGZ7k9bNp2rCqzWbyYReD1YMulrBCN9ku6YpGSPkdNz
KDU2JMmyyrzCA8JzAHrMUTRBzj0N0NO8OFd9USbGqfcE4QOvwW/NXbcetnjZYp8C
YA2Eu01+VyXx6kzbi9ARIa594Vz3OvG3Mt91aBsPUSHmy9F03H914w05yfNWSvEa
2Iw153K5dnCehMm/x/AEzyR4i0Sxg6Klm2GHhY9pFy3lkNBmR37TCRMoju+zghC8
IIynkKd4JlDk6U2KzgfNjty0pxyTq2HFOWoK12u2EF1NGsvl+lfOKg4JeOS07W7i
jveLgMduXm5N/6mS+0EQULn60Xmk1uCfJrkuoJMLnmw9DskrSTeM5kbDE2TECboB
1ekgrpVopMUu6044ep9VsevmSE4jZogMCVY5hid9oTcCx6MorNVH1qOU1dZdBQaD
rGznDv9Qj1XCiB/YPGcThcOVXtnnyz95IddBEeCSJtKDC9Xkl9rIUNHLV/nLL6vn
dgTFZXIERByIkyZ6Q7yqWSJP6bD7tkHryIP55mJuW+mTo/tQL8TEe9YhqizfxvGZ
hQpPTsgKpEi4MjEZ6t3e/V8u+tl7dYUGiZNsTsQqDxdXDt910mgZoOCZrBQvNtYY
Is8Xjkf+nxB1jYIFd1YjhGsYiYK5KO9P9IjZBgtxmNA=
`pragma protect end_protected
