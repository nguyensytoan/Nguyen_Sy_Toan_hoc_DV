
module debug_soml (
	source,
	probe);	

	output	[31:0]	source;
	input	[31:0]	probe;
endmodule
