// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:32:03 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rRwQNch5HZjp6jTYQTO/yAus09EHrc4J88TPapkqMYeL1XdJfXTswPfNk9LiWJ/T
c3YRBoLZtFJQO59u+iSbTN9DbDDrZCBd9naMfHmCr1n7slRHUnTXhPxderDvtur9
EDcno9XgB7ykJFCvz7srS88xQ9bwDwAJXPTOc7/B6kI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30112)
x3idSoL3Rn4B7nk4gLwTOhxUXhRsT1uCqbIo/W8zCScseV/y8ocKrV16Fl0qbCGJ
UcU3I6oZpfHZ/ribW/VFZzCdTi6IAgsiQAyIctR1CChaQbmJIqWzhUN6IwokEa4z
aWQvt6jlUdgOHgY+cg66i+pS1qu5LfzUPnaCdgxLlbJDTxx39oBbMvmSfOPeXIsW
dQDNiqpsJIsZ4FvJ6gb59M/JxKaG4lD0PaS18M+Q618YIAhrKOhN2fBTalnF0aN2
sPuKPzp60bkjXayqCk20kJdC9kC19Y2CmcvYSrEPwT0Tt1OSpbZQOll1o6lPLRtk
qK9TnTdvCrRnAc7YL2FmUFquwtdb5RQOddEiIAaJWrSTGCr75O4vDrjmCxqFzDgY
S7MgH7g6BX0WIGLCfT39Mkqtz5f7ezBu3pSovQbLfJt485NMCwQLWrLm9Bu4FMBz
sQmYPSWIbX7Pwye6HmqOX4xbCbiv1bVZ507qThOvt4Y6r5ynVcixqalpyUZWsrSX
OdzeK5UP4e2XPLlbp59M2u1BTvk14Bk0zyqhsi/6ZIhpT/0QmMXottbbhoxFWOWh
fDMU5P8edqH3Tph0p0sOU9ZSAfcWa9jpEYMDEkImdSZuIAo8wfJQjZRvg9yi/IzN
kn+66puuvj4I4BOuXUJqJdJ1E9GI4VA+/ZnW+iegXjJeEtG7+DNSVXLugJ4jPYsy
AfB2dKLkVyriaEQSW14gxueKirG9CcyFBJmakIEG3ZfZppC4+rIFYj+NIfijwh/C
PYtvjzlpyRd0TfUC5HYr8qjjTQOJiFeiuEmDCVlrD7svjeNB4kILzLuqe11L4aya
L8UkFvHWFtO2gjIPkMBvbeyMaEG9riCl//6/JC2oZakTBl9UK/bLc8/yeJraTT+s
3IML2A1c/uUWmSYfve4OfU4NNOsmoTz78AUWhvtJ6AlHi3PuvWaDTq8nUX+MexNG
3S91juxsKuK0HDxTbDh5oG8ug0mU5+8o/7f0Dl5gs8kcXYp4C3gcXpVkQtrte+I1
y30QF9hvHkAAilRqBqUz8eaPNOixrmnb8t4gT8dczdXERu3Pm9ChTqW8pRgSfR0d
7A3I/4HY89DcBjSkc+BNv0zeyr3mnL2y0mq1eCJsdpzXVbWju+euo+Wm/DzKdKJI
vXRcf74oLKsVnqUg614r79SSbVAUorRMmty0N5f68VNvM2ILWy+PQFvhSy4IbpyD
6p55Bj9THyagasaKisRiUKItYkGb3yMdo39zrGPGF2YFcOvKFdZG1hOBQVrAyfRL
0JgNC2TN1oQXpJ3ARS4g6UNB4cnY+4+TUO4T7bLKvwYN68AGQUGlZpC9WQ+0mmcL
0ER0FqHn4AWNZrg5AuEfO1sl6jp5259+mOVGhdUNmcJekxZPf+6qvWXCQWkpUmJu
qZTaNNcgIu6+hXJXgzsza0Ka20eR/78RvyxW4cIcwdwM1hAYFqpIqRNg4kxvkQB3
Pb4COf5Lw8zW2aaoSrSrvl4zZ9GYLsmDHmrezdNEVs9ekEQDRcR6O1xzHpe1cX5t
52x8DVmBnfz4jlIKI7ndpI17I+9Qn1/Pys/uDgicnNpRIbV7d9ZENXruvxUyKE2W
vkYpMiW+lFY9RxIv29Wsr0aiRbo1SO211UymlJLOn0hGSzd/Hi8ltDJug8f7WcoT
tix/tvnvR615OC+MSbqh9aQNPu7bl5NBlMKWboXFlxpUq+Vq2WL/q2us6U95GzsD
0jecGU9201fV/tbMMXiLT+gLwcci3p8WkCyXKlM0ogbwkb58OWk9BIk93RAdPsa9
gC0tZnzNBD++CH60uJecniBgJdqs1GZdX3yQ37NowzGhlplnCcWXPTs3lnBIMnmr
nqy+qcUy1uxSnB4wQTjL3V8A7m7pixOslRoxJisGwVcClX4/r5yG8LYmhOoBFjeE
gt4h7Kn6HxRrFL0hwoSrz65zYB8ebraTqeDpsUnu0h++s2oYdjEQsKEursp28sS4
ZIARevi+a3/nSL7XJIxfAfg5AvoS1rtjwcOAAI26D26wygMNHnYE/YUVMlK0Feyq
C+Yns3pLuONcCZehnd7E7RGbKl832XEVRaqLl6xgiOE6zZjxYQlwDJwqEsE2mImU
F5hAzEciS8d4O1ZTMdoo1nC9KIcZflY12ZAH2OnKS7ijMIydH+lft5XS58us6M1m
om8JnH3cG28Nmzwpmv2Ug8cyNNcSCN4tiOoURQRl9zIjTbIAtrTT+BEe0VAfbHfW
PaN6JrajgRDDxwlpt7DWoKGKJHw1qAQIE87sEpBwTLtCyAUqam2lu3H6yx15eIP8
pwjFiXTK1r26zuSUcE5J5qjSTiPrcbu2gaujMcW53T1U5m/oiWAGiY88ZFwNcch+
V/oO2E7dwkljsjH6fJdgPRQVqnmop/qqn8sFk4pkAvxCIghcH5jHRo2iHweVteW+
tKanfn/k2kGzcrESITseDNWD3YOVC9kS3UEFJ3VZ4CHBTMuii1Dqo/O7pVE7x9oQ
W40eh3e6odB3OhdczoL4oUi0T2J+B06iDtuJAZDPE/mVnQO0OdnV7dqPQTdoNEGq
ctKAuOIjXcCwleOIEtWZWVzow21YRiPws6C4fnSt5UMntVdw1c9ygmupIF+VxgE0
VbJUeBMDRni+zKo+Wzy/uVA4enEsj5TYCjC5zd0zT4LKu7JULA2sWJkFxtzwZlbn
fonObnla1sWAR7SBtSsRGD4gUGL4wVHwE3KzKSfs4G4GljszRha1I3+xyM4OI/si
1uZEZLu14H6WSvkeJOj5/wrELXV8vDCyDdLsYfJe1ikTdIYmmeSrjzKo642UDdeQ
Lykjb6za0rhGu+ca9wfktpZbCnJ7GAFtiPe+2VSwdPIM1/HpzZJ6Ea5R5yZaB1UE
f1x+W88eTzEg4nWyiVb0BQ2c2TkW/GJj5IwxLxmQEkesocxqcEXjw4bsKopRswhb
B6SjOZt/jPj1iWncwhfp910Qi372/vhHlpfYRWp/yCBmZTIWX9xWi+HYiJm7zAve
3Ie6KOUHKy6jyWBHFLjBdFDSTu0I2qPzPrk7sOVER/SDVFYgxAnjoGhlsoBJuD1f
TLdetgrMSr0GL8WL9xyCkjpPj2GW92DuGJzXv5BFNWjaLpYjSxnzk0tXQY6ZOBmc
cfdY51RLX2seTr7OFKMOx2AL+NPGTLB3kQLPIs8P7RNG2lBrucsNpIhEKkHkKJJ5
i0JTlWKq1P75Rf+SFP2T4u4SUVDOQPbpVyBxah5QNSTT3Pv3jbd5ogxCvXtT7MvX
NVchMfQ6WF5O3kaPqvbRAIhOyTfqE4PFtZ033kBXHm4+++yQBO3ymGq8Eae4Nx9Z
PBlj3gI6KXMuanV85CNQ7YOFNQXi6boFA2VT3vPbOK7aiLfXYbf0bDREAjqwdCAr
r6o2qeCB8PEaeidg8wKVkLpYYRimQIexQvds6vaQHPRBKxAE3SjhePjQMV5CCAGj
Isr0dI5rsBpl0EWfw/SdYlyVZ69O0obpZLNTO5Lxc4gGPAGCAhaUp/Rb6MKM1RYm
/6zi6yILzH40M+OZ+qOo4TAajV5/iGjPcT/uxM+j+3SDJ+iVa5ceWZj1iiZSuPif
KuDWv/Ik64hNRfB24bna8q0ZTVxsDcnmSkrISnLPleE9CFbBS+A2d6CCFI6dAG0S
2Be3C6pMKph5wmFjC1jMSK/IG081fGrK67aOxmf4UbHxmIymx7ynYph8VWeKnuYH
QgxmPvLJVkHFGNSVD40F+n0h9pXrVcfboDYIN/XVZMKJz646OIeSKh+J8vTGqYLP
1d0LgIlO1VExME87Jve2wBau4u++4SFwFnUV7g4Bkd2QRgOIH5f7KGucQ8rEoiZM
OKA2IVE6sa2EhN9ukzPAp31hUHNMow7sF1u5kwRk5djBTu2FE8NfOxoSRuyD9jCD
Zw8H/UIYQgbiPzarlwlCd6F4ux8fbVCNyenPsY9PR477Vl9m6qlGPaHndiUfDi3p
N8XNmBW5A5TtMV0xY27xZb3GKQye7c5vWjddorgz26FY1GgJSCdIytLuQ2FUhWYb
xkCi211jtdJCjN3zFq8k0HrOlsD6Qq6aJFDdfxKbfWUMwSeexA5ZJQaWBhDSjQHE
U5kTI4w0hIHonxq2yHSwkHxpOOEA1mv1gG/0o/ASucAxvdJAwPoStl4p3Yns20N+
XuUKO7Vcb9fsb3VS7DBcAdFhWmLF0cdmhx03hfqbR1jn/e5ObULDXSCwGzc9MrMl
rrq/AVl9mIsXSUkRxSlej7v5pQKld08arbnRTEYzQKuOH6OwQkNtbatLAfKb9vtN
BMc+JOayfaEgYCqEEcGXIAmz1+Z6hBrR7acHb9rVnhfFdZ2gmMGQenO4Op1yVvIr
VCkFoPw4Elbxb4ZdMCu6Gi38ibJ8kYEKE5ixejGyCUbeAKVh0w/q430XBxHKmaxg
q+PHPHy7aSrXJKxhj/48d7j1WH7VdWWntGcRkIitKYs2usGsvqT3MpWagkMO5pcP
ai8RM6bJzKdaYTGSYGaFQV3ePr/qUTM6A9O5FTkIeG2acIFHIz1J8ugbGvKrjDDB
OBypB6qRf7EQ8W5SKUHUxRSW9trSCZSjsayR4ZQI/tb8GtS71x0DJk7fWpIMztp6
Wv1FrrgNMrQfr/tbKjDST4atuJhzZfYenNUmlNRZl23RsK8C41FZTUCcrOrgDz35
YqpKt1JqeQMEmFBVy4v5ZcWdnhIx1Kxzr1F8qdueczOw6IZh73h3FIwIumOYGMH7
BDvDH3dAObypq+5YwOT5nKa5BDDSTvhaqmSJf9avq3CXc3vrqZPSxDKQTmELvAWm
hfGrBm3VtRe88upaAEtt+NQKXp0KFzYH/SnrPZ7TUDDKtvS8kZSDTpUBBhhpkxUL
+S/d/kNQaIRPKeKFOnSnBHBn6sNsCyNyhHVMvA90w4k10pp4V0bfX92nudp2XtOO
zCgsaDRxb4POmfZDhGwbFCyA5mVnxNGuPaYZKKPhFCYv0pVIjfHOrnF7Ee8e81q0
UBB15yOe8JDnE0hmQC2lqVvYbhkRywa97IXX+tzdjWbyyr+cpfrXhm3sxokG+Q40
OTLne+l0xM65KmI7MMoG+2huHhmp4aXFK0DzY5J9GSmIlcHaWEogqwarqBIuka57
dCmo/e8sgpAsV6Ea6ufPesP4VBfSE1EDMFZBSXZ68P4KCg9msNDSkO+T1Pj+eKmC
mMzgUeAKy1utLW3KRfyRV1/HzTadOBuiPdDhQnc8YSPPUoUzTLQ9Wqzertjwydx3
HcCZ7ql7OlCn+wmLRVuOIwVuKN4tR6/ucCJ5NuFdksxzZZIxu9xF7P+gUQIztQCL
6F8bVg8p1UxdQfWb9ykW5+JpcaFOQOHnm66UboyIimHqPLrg9MsM/6rKaSmb+RHr
ugXypuOXLwst48SMpVnX32GqnAmo9KteDt5pX+3O3JpyNhjO6+6/bXiEzVQj3N7z
fXyNPwpnFaLPCtRJIdII2T4CxmtZ31y69fbBHmP2VhFP8N8vjJ/SQZbY6SCz3ghH
H7SyhF4bwKXHBtX1umE6JZAkehw4TR/708RSyk+hZQqjA4+l4lNRKmzePg4WD7i3
6fDCkEKqDCDzUEugIwhudru2SQiO77+RBHESGktHJoZ12RaBBOw/8d8Jizn3I2y3
ROkYNaFawEC8gexDqXGfUr2N9srMWZyYFH1i7jT83KT++boq6aAsryAD2K4hMUjV
0Wlm/lle5cNPwFAAPP4Yptb4pXlmeBFZ2FCUBsBYOVBi9mOP+0WJv47HC8XgWnnZ
JX4v205edxk+vZpXHlMUUQbcVmg3BD8/Kgqmg8upG0+rrWSOK6KwHmfYgDm1EQ4M
pRaXtoMXqOO5wff5nYvteMf4/FIHDaMuNkkK89X4dLNJv98BR3nPu1HoZ9GGj95B
slaccA2ArW31uMDslIzqJ7G5FY1/QoQ+kG+UX7YC6GRlcOvX7+81+76Z9uy7spLW
fqH1Q/kvjtLijWDS3ACdm9xSMsg49cVhtf5lCBB/apQ0sdchWRUoP+tOkdgW3LC3
qWDU907ieovzHG2aIPMx9ydmqml6KFWBNF/n8hyv+pmZ/2R1gpZUqu5ADEZ0Yv6D
+DWZHID193CKxbpQaV/9FydstDzqH74OkH0jHqtTKKwhopQ/Y2gU1pfQuQuMrbzE
PZVboaVPb5pjRB+YfQzf/fIoyWpxz8No0QKgW0AcJmnw5ndRHLjLOwWn8PHpBlu3
ZM2edylkoN8AyqOBpsZ94R5opC3BF2ctouPKqgEosxOXn04kYjnXQ/Y5LAlQm8ZO
xo5RcMGV9hh9T+pG2ARV9G0732qBAvcFXzxvAoibbm/791096sxHfP754M8wtJz/
4jWA5egPwc8GJ+qGWv63UEOB2qdqZEZvGoPMLRIM1ZI8NJgEKrWKha6DM2AWXJKn
+O64TByvG4bbk+ZXpafyBDaKufoj/jof07PhuN7TOvnBHkvLG5jxpghnFjSKK9OD
9WLscFpC1GfzldarxrkL54XL4PqVIOxwnK5a1R0hQcseFhD2uF2xMXj9gDKje1AC
yTK3AgVNRzjATLu1mFnLnVRKguF97i4wJuGkWBhi1Kh12pHnjL8iDK03ZNBifMpl
/Fi4A/9Sk846J22c2De0KUnJtWduhqCDHzKgfVoDU0JkSW2r6v3t43KUj4PbdABg
2ZNjHRvBBnTcEvvQ0BQsq43GN35PQ3zjT7NASsqfuCjA8cLWBqzgoYgWUSFlG28M
9mOThKzqq6f0gVOLuQ+3TPJ+VYfJZgsIz01quZ4T91sezHKET9u//5VHcySZwtY4
NS7zR4e3xLk/McPpFcqEDFRtHPdxVjniKlt8Gl6Ezc2Ry0p+7S8kcYm4U+IPiqKE
e+A14lLXjkt7J100J06c+0wGOOBzdtDOWVdDRPtMJ2yzEp5ljBTnnCFG/qcE8oHR
EmXmD0T9dbdQ13Me+62AvpRK8O7yDaOVtEScB7c0e1CCahstQjjlReJ9e3aIBWvq
nJoAjUUAtDZeEcBMBW8lqqJb+2KDP0yV9C+SgU8IvZmxxA+pUxU9kmDJZ+ByH3qJ
ODZ9HLqSDZaIVrnoMxa0P9VoNQu3iuaEpj92ALaI966KJ/vYmWRNjp9OXOeL/H3q
U2hQ85O88kuqdncOtOAxGoogA+V3x089SMWInbDsqoJTApZ/R5NgfH1apwu3ucyp
aQjhsp7iLDNE3fXSGgjyziOcB4pwGo+5FRuKoUtOD3LLZn8V1rr2fnheAbd3m1R5
3b6PdHAgxT220k47/xS2n3yKvbXjxVaWN/yMZ08TxUI+gmQznGa5zdIuI6Ro0fYB
x0/KPkIo0p0ujUtTaWCpPRqadIuWLTkTi4nbkTQw0Mojsbs6Pcz6IwsuQacbQNKc
wdiUKTnT5otkvyo5McU3wXHKXu6DLruCAJJQcrvfH9ipvemi3uE5q5WuRxM1W/oE
QSNcAAlI9UNowbMzxb3FMzSMxpJN6vxQlgEkLuUDKRDaRgA5G6GBYk6GdRYxmri6
o/AbaC9qqT0giHWe6F8QJxE4898pqaehGoL8zwzPyquJal9v6DreviWtsQeGPux7
e6Cywtc351pQivl78D7asRz9GvbLOpMr9dY3hhsG5q2k9fhepEJNzfIddgtnVjRQ
4Frj6gxhYawUtG/nCcM4AXjNIHXb1+6IfKYUGzZz0MYWVfPMGWFjFEMQne7e4C1W
Rg3LMp4IIn/dRFq8uL8ZB0bqnUbXuauQGGbFu9jar6SWYE/+pYnLoTcCwQo5cZQu
hHJEnUi5tts92FUFpe3cz7g6ck35lXcOo7x1gWcAnekUMXlCWLOalcFSrWE/4yc5
sqNANcmzFqcUa6FLGYHSWDf2AkTiR2uAnBEr1hDDyDPgRFBxff/uZdVJJc9nnaQl
G64j+LtBSsKOjFqZqCj+iuzQ/qJvg1w38P+utAY00xRiJVUr4fdRRvILySP6SSeX
Pl19Mx3AGWdKsvRYGNzY5IdY/VEMTsuhsQmproUjyObWdHga+NDOAdMUq93iFXyU
rbLl7zd0UpFssKm/EAZJQeqHUN6Siz3HRxJ6deb5D18LliIB8J0Fxam8Mk/awiQ4
rKFZWYmeFyGf5+HzbVS8V+e3a+8OJ+bID+vze6+X4Fq6KVcVqHrSZjDNgsy3YPch
O4ynSM2W68Vzt13hfn3CY6ihvMxCm+ZZhtHVh6EWyo/T5qXYzxrPMWJORIXTLqup
Pa4mUhrJ8owKsaZ7l7E9fdu8Vi6ZqTndh57nqHhSWK571orPVd0kF2hgNQEhjkI/
qu4Q51GLOw7CzD6kzTPNUg12vaTJnlOmlxeSUd+46agKtj2LpqVOUGxef7vVfcYv
xDwyDI6fGGXPy4qebptus+IXSSB9aRrTL1pn9DxI2jr3DErS07iV7k84rZcYaBIF
Lsqt0iaqDziZNk7vdeHtD/bVCs6YNVYKNzOv/Mj7FfzsQTpU7SIpeN4K/jKkQUG+
Iv756LxYfakX/Aa7dII/EYgxfOIchevBDtfsfvyqtn1xNOltyH0g7l5n3dX4b4HN
Hs1PlTWS0ORZbdg/BOSe0JXaNOlWn3o5eQAmMAaR9+5+kjg2t5h0bvnmTwvL5aZ1
hDRm+zKHD/uIw7ct59IGgePo/VqsjSgThVg+DMa/UqOzoPMz4xmHqzbTQZ+EXndU
Gt1lbIYxqwjvovoS6PVbElkcHLgPwAVXP6zzaCIcvEe9L/ZVy7CPiAZO57xWNQvC
a/uB4pk/25P40pboxWz1CKWHaeCavy1Hnfu1+6hMJKBcAxIpt0W7TAFIzQTR2Oj5
x6DlgkDLM62Au5O3foLB24qO38c6lc8YvgE9amalc2GdWZMGtSXINiLyHvOfmMBQ
UupUaE439a/1uBv5zIAHacdJ16qhXM+cnLOfz4l8pS/A2R8WWYTy4/yQAZQeYQWl
ctTLktWrn8ll9NLtqS3HAbBD5oeLnnaYg+JTY/nUNSdGaQKK4sct7tCaOaxZ/BPs
RhldsKJ21ZRZBx59CrmGd8tIdnkWmrFwpOadCCTjq/k36HmgUNtpvXl9NS7GUQzl
wrI6krURvzQSOTEu/H5T9acRRoENQ3eCEEEIe/zpAhTP/SjwVY/6wtpW0GF/G8DS
d0yExpbh+p6diPpjuKsYcB7ztWnaP5yT1cykz6AJ2he8xOPjrLfArLhKkQzTKvs+
FlVKADRHOhH4briSgaM4DZ91KFQ7Xe4M4clX5hDsCBMF5HZWBAnu7ElrvBNDkUks
77bwRGZN1MP+E1f9hSDPM+rba+YDWsxBX7HQpyYLiWzIdFXLslln3o87hveIpR7z
rGiq2m6lVZpj0BC0Anng/iL9f/0FcspYmB2mK7z9KYT4TYeadM2UzWmGe6pPtJ+h
ZvSOwluMb61p9nPqMxhE+jUSK4NxI3qoH1Sgu+/6snTlGITo6xJpmEh8l0saBUVi
ySjX4OBhWOnC9YYMxj/p9/BcQv2h4JqFrPJkuL7hUR6IckW45E2XJ75LZSLizN6R
3E9nhHmpUSbQfY0nQ+lfHIR0KyVp3qOU8rS0Bx23hnJCUN8CbNmc69SDqkNDWcQ0
b5zPagoWy5CoSVxTV2/UNOaKwb9OwGvwsAxINRn99D4WLs4bevEpti+7qou2p/ki
6WF/DE81MsNB8SbgSS8id6DSADa+F0mng4hY3ehGNfr9cuEN/RySoYuha+0bz01h
XTT0WMVhyPdaDYZXvTIfRdWT6SkIQneEP7L6QyNWbkdXefUY1D2EETb4c6eIDS6k
RrZ7omwgaI+DQPi2Cp66Nxh+btkq1ufTU60MBeLXBtoRb/KLCaswp4rMW6SoQqWo
XB5bpDc9VZ2EQgJYzcG7TDH57H3mYxBu4R/gOVFUb0j7gT3Mu3kko8m0FMpRo5sP
6YEXF9tlwY5LDnwhkNdDDdKIHyLkLBviqeWJe8vGzExk+dKhjOjLF3I7PUtoHXqS
ChDyESAjhVyI0rQZsIpnUFOmady5JGAnWv7uY8lo7DBxGfe7tVoLGlZTkBdmXOpg
T5ze6kre8a+AuwORcQpCbYsxTQ0jOmGFbebnXFCzaITemTYXPZIWBs+41bOsxk9K
i+51D0ngwaDz/bpIlDQaCqqIk67GmYZseAX5O3/0qX+f+x3smgczGqlcIsCq+BE8
sdyHQidmsMNglH3Zgo9El+JFeqtGNU9yx3tPR6ym1wW+Q8nOEPbmzea/fHk9noEA
Opoj6ayNQXl/bZEAEn9ONYur+g2Dc+APicRubrT4nsLUDEwiMtHTPvvLmOf4cJCq
fuI+D9GA5hOw6spisklZcScz0JxEstjiv+eu2zA6DfHswhWku5kUUqbt0h97HvrP
O51CkwwfUfqK281K9udm59aaAGRDQemM5EEs2PqnQe7tCVPzOqKo2rijqFdIlXx3
oJaHXNyhDKogArZeAduBEeZfPNnIgGY1/q6Zz93g6jMvO9PiEq9xKH0hDdYBZzXm
kiYqirtnjjhZZ1J/x9hsBoSHRaYPHab61FdGykjnT9BNzcDbE0H+RMB1DFKz2JxQ
FjPpopNNdQnUE45vHNWlSlJB578FTFRcM5HCJYuy6MHFcSryGe/585ghJLsehp0p
d/uQmnLXMPBpn1FAgVbeB4yOc5CcAVYeYnUudOsMgpX4ZOmoHjbgb64CPWa4HR2K
Bfo2HXRuFl8/JNJuHbBp4KhHvv9Ww4ubfo7IUd/lXC86v92NiMoLT+wEPGMZYcxD
6+dM4XqkPi8Xl6ErJtaN8HTURgGdkiGV38xxp7bR4rcSaYcTFkKpECnIrmsGH1K4
Lq4R0DzuO9bVQdLAzroOmG6OdqREFd4y94z0EOOHu0Y74hGRa6QeY7gnTI4jCeyv
c4nLBeUmbcsmoRI7ZvYKP/4Wb0RRjQJ2rgRQDniiUQxqTEhqPht7pmS3M8FkWWuK
PWPHUVe/Cu1Qkpqp0kT0qpct0cJwczDX8Etgc+4AiWuc/CMlWiJjfj4hu3GsaaOn
8bELq6XXPTJN2f4yljuMQWgM7GzaiFNi9OgwI/ingwl9kuF6GFjNxBbbTW3w4QRw
JSsl/z1e9+S9w9zjq+/BGNrD9zFzXRnpOdxd9BSHgevkdXaHeVxlInjKZ0Icjd8Q
QK2K77SWDQz7WMz31SgPQLzK/lnFirHspOW5tkQ1gYzs8BZ8hzxJ+ubX9QfATcek
ObxSDt83OcgI3LeLwgbjV7g9FXJ+V9uVjOlGq3K7mbGquG8MpgrCKth/HnpBbpOU
TTCxSbxPrOw8IYvDb8xiZxnjTDxnan6yv+9rKYGMEDis8jdLVzimImX9szTAanLS
hQbUj/MkiCmYgY63TRHstAiO1oPuBx0eg9JBojyiNNKoVz8fq2nEOcuX1V+PzqaE
BkXSIaLppjRfyRdX13iIpLnhDYYhNHkDESnW8/vAClT2S/rqndl2bh2OmWZAiaJU
J13f2sfskKSpjUt1n+2H4sdSGeakAlQSSdsVCfLeRI7PF70Qc/rfQRXdgeMVZoOq
R0CmjgTbyl8JyVVbNqfljVWvbO4b/d8MHYevon4ti9q/rtBjWKJkejgGv+o4LkJ3
pDWQSeArILbvHVaqZYb7fDFcbc4fh1GG6XOy5m/TuGshOxQSe8+DjBRqeVOk58AH
5Z/ID7pdeDpgKJN9D8EtE+NXa+WyQFVtLR0+y5n/EqazBLwhF7n8B7spyadM2QMH
92p5THksw2dKuAeji2ZcswykgxL9jbDRb6Mycg0oPoAOKqhTYCpMBW/00rlwJDtp
4SX6wPWlhYZMJCcj2mF8ctSRaa2LWV1N7yrkzWGQU/rx7rZ8glToTahEGbK6HFfd
lbNNOwWlTcYtJMsED/gjXgbrekVInNNapRr5at/du4BVW7q0jfBC18M+ivAzHvH6
DyNKjtaLFCDOBlTudzZsXd+hryHNQ/I8ln5Ne5U9/PhPcYWYtMr+Q0YO7r4WWJmJ
8qyAWHrdYSjGBpzbJOYFF4t7OPFhKDUovLi+xyrkKEscpHq/H16JJZFABytH/Yc1
5+sUCcQfuQ9k8xx9Yzogpr8WkAShH6txrBf0hQRa1a+9sI4tB3py4ssPwfWPCD4F
mYGX7BGxg7XeZ79vaX9Tu25Wokf4tw1FZkV7iF2Bp1dFdv9vBIYIpvkpRB4sRHYD
HiIZ3pXTfWsdEXZrNmsR6DlyjthW3XbfiDHmpaMEehT9dmktITPUA750/+KsIWOQ
KtxhAp7NY1rjVVTBkz4sbJpa8A30jlp686ihS9zAy3oFJijdNpbYBzs1Fi3/7Ew7
rRbbnM2Q7GR6dcuiJ3zt6iNIyneyVL+PJ3sEXqqTT44xouzYXJ7eAV4UvIn+MOJv
GLET8+mhAqp4xZoG8g0GectYhS6izpPcS4FyYI8AAW/6jsznQSMzQYyuovg0mps8
hftn3mSatP+8i76/YBgoJe0l2mfumN6Vf2jaAu6CU0CS4omnwV98AXrWnZI5L4+E
uSIsfiCWcl6C4TABZyLRz0QmFNeOZz2p9w9/zhIhsdMAiMrHpEozfzUXgnsrWOvd
pK1b6/0cL6SiQoqUAFY96uz36kvVj6BUGoSLzeotNJJnk9WEzxqzS2M/uXZPPBL/
osvydyEbzIM5xSKoCxg1vsqRAcNqIaMr9KfCUOMVeyf7lWPqvh8/uYBbCPOiioO3
IR3EvP+7DSnPG464aT1y43A/zzS7BlOgfAs6jLIOGva8hZDohi7M8VFFGioNlojC
/95BKoS5RECU4mAcaOqF757aIOgtyKxX5EsjyKD9Heccsv093yKECW1X/ou7kc7D
VjaARr/vjFf528P1TdxIYjrvlSOETaSnZrw5VrwcKbDfJIaBBcokCfwfXTFUp74x
t8MJIwGNYq1+pN/77W5EvzE+WZ+WIo+Vj/J4amGz19pvGSV8Lbb4vOAhGIDRUB3T
UzuD28S8RdhDCHxdkkeM7s5dOe0IlHkVQBwcAw+lVkoeZ2cFWTDg53lnHiqs7Kbi
jpXHHeor5NQiVSsj9KRvXsTVDLD8IFE26Wcz5/9fq2YXioxn9Ff892FHFTKKBV8x
YPh39GBxLL+Uk2w4P+B+XsO5xggoSE2LWQJ9QGxeB4C5l8b7fj8Tai1BnP4hQ93S
ojOL0ZZLQw417V4Sob9PAY+vjjqc+f2KqCpaKM7IgjlJN41gZdDnaxSg6M/W4Yft
EEW/L9SCLubyxk5SPR6qIyzczPEhu3DwvusuGj4QCM0ze7rNFTaSifgJmx3om4xq
2e5uL6ChW/GvfI8agskq8BMTyXoM2g4Dqg1yc3IlS3vVaDTG6oI1twlcFseEB3p2
3h3E7Aa+CQM8lMXwUK0HgINsE2u6UZ6NyzcWE3LqpCC5XEsuw4LUGW57paApQmkV
75lZWMGe7w3sgrfooyek66oB67WIi31Qyh25LBPjmszmFdwmsp7EcAlJKERlGcv0
YDePp2vF894tSvUN1BwUWbizAiFPG1th0nBO0QIX+ExLUS2R0H2VBdGm16ioJB3r
jeBslRTuStz164DJl8BBPA4thP6adQXABaYoFjhJkXdGtMvhjnQEbSUHNu63ckaQ
Zydpnzr7n0CtycUc+jpl9iCiuK9TFBtQB6a/IWyzmCowNYK2rQPRjstajoFBv0e0
BkrUZ0ZzYmae3eu2VULDe4GYSs7jnEPzVBoLiFh/q2p11o9AYLyCz3EBHpwyH/2v
R63xjFa2BVJnBrGh4/d1AVB9V1LrzCgdv0m7HRGkBd3XvuRvfo5CIa9/v+8bf6M3
ObUrP3mQfdmup5bMo3Bl5+6GLM9WTsIXa5cZdJzzKBaiZUIoWDZJ5vUuzzdI73V2
g5tG28C7vq4EJI2vRQeJF970JfGFxoBH75A1j7Sj3QGU+Bp8KWica8xAkfzrbQk9
Zeelh3pIbAtXnATlV4/2cjIc50ekVc8gpiG+JYnYPXMZhdqkRw87o2Oh7ij6ppsO
pNOrXMGicifCDzC9Nknbnvd8X/s3PlMFYf4XTVryCijULhcGt7a4sKgYya+AGRSi
KKL5bKfBYjIq6FU7jNn41VpOLLrqk4iaM+y038FWFujEpY2srQhpWC3JM31GaAzL
kB8HJbMyDpc/9rWl+OXuRZZX+MB9fDdtyfl8xZW6lGBJOLVXgMMy2IrtBIooWZRf
TI44j32arPVeNAMSsthAs20LHCZuOBtEps0/795dKCs8kEH8WEWMZmNnaeQv+Rge
WXTykun8UqdQmNhU22mdAJgFP4exddk4yNaJD4zqlv6317KVfNn2IVXrSng2SwjU
i2ni2Daan+yZV0i7OgLBHGvT4J9/jYXLxqhq44FW8Mp+cFi7CxEksELZTiRbOiY8
dno2+onkjTcjHaTtg6BQaj+OImefUb857xOljrT5WVFj/bMq8xhixIaFnHq/JT1H
c3v7SrzC7T8yWVwJ3QfyFgWLZduJxBNG/RINc/Mn6qoJXhBiHBoBwCHdFhENOWpu
Eeg8us5r4MGZr3IL4F4eOZIH3FdQjO7ZwwPWkW8QZLZU6go9/jcb9jDj0G6v9jvj
nDQPdu7gY/FVckaTvQ2W5KrP9ElTT7EOeJvYVPjTbR7L6YvRlHgEusS8aNbMR35/
CoricLXLJyt+bUgvYP9NZRQpSNpGc45ESshk5bSIee32lSEzykHBha04vRrFX50M
kkfukFu3fLXjam4mGcxGCsdKrCnvvGL3pVQCX1GDxcSxz5FX2XJZkOH24agD09bi
k3GMIvl+DNKcvrVKwSVcTYFr9xoPbLHcESU8FwitmfkZUMSt3gINkZjbkom/iUlF
lGyviK09LJgn61I5EPYt8nPHMciAjblAPA6Pw3mytd6HUu4SA+WLAMuTYiJKzBmf
q+wR/MSYn5IRWx0Y8MaE+qWdOZvUWAdHIq1CT2J3M0ZV2RhLlNCb4zmxCcyUq5Lj
qfWR380VIWNtsCBleZQ0ZEdf5wvOpVrVlK8LBn9tOCOe/4DyX5AeEX22d9ffyi/P
V5uCZfSHjqCzoxxuya+CxFvEEWBxbkX2VElXGWDZQ5VTW9VhTrwgXiP0yFYtzIng
5KsFOSYwTutnM616GAqoHlVXxC2T0N2u+Em7I+qCGOooU4eANaJmQ+VfWHOcO8WM
dc4WrCJzVKXrHFMWLdsCGpKTba0hZP+nQXgy2jlnw8UmpOjm/uumM9bDEBnwkTih
PwCzLZp2cTC7GsGtvF3RLAw4qYXGY0kZCbmqokKN8S4LRqMbWipnzGGIx92xWvYN
QbQMJnGrtFhK87ny72lGNVjcNKjIjxKgUm9A6Etvb6I4T2jOsP7ggmXlv3P6JL62
2v+jYVMRvyQDGo93IHrjICXInDMLBLwXMXzgTFQb4ZRFdIobjWG05bvluyC6+h3a
x1kl+bZOftflWVPrwdWFISlCnDg09li1AQiPGDvfMxMUyfjeSD8NWUUSoMILn9Dx
fHd4Hm3Z4O0BuEhUoJn0tOaOVofSKD/YnvktcKXbvDmA4EgBdlmsv29yH/VS2q7u
roYQQb8Duv8rjhmlHriJgMGKPzPBzgt9Htpz3eBOfpcXqq9yKJx8Yf7fnhy2vJNs
Z3fIwcyaNpYTTFscpfpGGWub8SM5tNsc9Es8AzNE1PBeg3ZmJuTDosxK1dVhZpK3
mxq2c36T1yKT2JaeZFxsBsRQXPfw/hH214hJ6QcZOM0+EWE2nSuG/kildbSCKk/n
LJRomaXIqI2MYkyzBgjHZe+Yl6OFACcCWtp59hTDnkbeacadCzIa/AY1R8RJjTNC
2tA9PlYSXO0RVFNHHajwQYjl80ISR0wJspQ7pIU5bVfvfpSfflpFu+WOAO5Oj/Xp
Xqlp0a5jxafdEtu4jp3tLsqXMVgZ8YgJiE+3wCG01UC40d6DA/+yBdgXK0apHHjx
cwiW2Wb6Qm2bb/0uV0aRNz3dvrA/1Ay8yWrBWIWIpq/d79Cbii1phbyTROR2NL0g
q4PJJGHS9ddj/EUiEGcsNSZQsE91Wcl74NBdMrMSggCIGqzDSOYzevDhxRoagUn7
oJaFmX+cBoC+X3PkHdLbjSh4Z8fuIW9Bl5TVancbNGULi9udH4R0KY4xe3vBQIQe
8NuK8T8KQQmpQnn6sMC+RJgk2nP9+Ib36j17XOwKl3A0L1S2XbU6EBY7QhwVuTfV
Ucf8Jfbn8fHBq9Ra1QkbIUYgmicbEwZDS8JsZ69YmJ/Kmt5KkMt83A0w8wPc3C+u
vlhoYm5UUDb1HNRAYoP44k6u0ZiFhT3o/cIynbd0M64vjHFDzkjs7cFQ25SyY/GZ
XhCa77gx4h33jh3tQfYoJaHrcv/w+uDgx9Hj+uotWIK1k77J3lgT9VG8Xq++of2J
V92/ULb0vCDq0ZiGg2iAN1eCAxVoFVfMCW/z7X22/epoSr/V8iwX+kZv1MTcQ+V6
0ycrR14VWJDzRI9jpd24eHhVnC31ZYI1ixKAsqaM/ZQ9LStmliqtuSFf+synzgn1
rtfJ9XErti4UfcLAT0dQnaOl0apJx+A2Lyr7u9pY+U/ypk2OAvv9joxMfVvnF/9V
XDLGkINFkZgb/VYb3pUG4rr6PHt5XYQuWRFhYBmjev7cLPwkA/rwz4z/tfVTUquC
IZVObqFechw5xvHOMjBkazZRUpTwgKc3dtrYTiJJtf739tnUdC0/MotXVbJcM/k3
dsn8s4lTEMhLy+KJen+4Y8ZUsV+kvpiUO3ap251SuqmuPHJ06T0fFUQ5LMaS0Xw5
k4n05VhVpXL0Fk59bbz/YSn4Oe9VZNl5xwB89TW2/0KiW3x7lxGa/0JwfgsNCpjk
hjhRxO0pYfN3kgJN4tWNhQ5ij2SkMOPgNEOu4WZLyM8STW+HiwX2PtTdCKfducQl
ccOcnHnA9KhsfO4QEcIixQDaFrgMPXH7XnfCKSTJnEvrpaVBAecIGeL2ivvLWz1A
dPb5cF74HxLOA42KsHuRKFEIfGTAXQgTQT3SD2zxtyf0v89Bn438sncNmqttp30t
IXotIbEBTKU0fkI+vUP7DHlQB3vA/Okd6ReeTzmMoAgyubGFDpmJyQRLlhKITRm0
j6F+cW45V1eMehJ88TlW9duJEodniwFeeIo2TyJBUWiEkv44A8ewWR3bi5PctrpS
UmDLZqNPRQHHAld7VsOt2OVlMxw6EKwLaJ2/njA2iHhMe/M2uw128ha4STprlXgL
s37RieLPROqHggqz8EAKh0F3PmfE94TVmiPm5j6IjcNoYT9lZ/hTbTQPQwrC8D/h
Lnms4XWWR8i6N7B2gp3Ut/xZ44oJ+nzHU7aq0HvTL4gh64GlOu/fIvUbHT1yTaBm
Jb43Eo6r2W5DD3OhZgZQmxqmSxxsXZwh3zQEXf336aC3vWoZgS+d7MlygM8r1Gq7
yVyzayx0VyF9uFTzuX4lIIjQaoQoKAwY8oomDqfyS+Rc4B6wY1YhM/haa9jEpy6e
pe58b/PCUzoOZhlPoZGfxuNqlFOBC/+JODd4GuVLABYogK1zIhzrSUMkCarIwY8Z
a1Wg5mGqbrj3UIeqwsG/BcThdhoxnUjJ9WI2eUKZ0C17IcF1Ve/FkDiKavB35K3b
jJz7BPILTd5VN7lWVHj56tF7RlYAkcbqiz+rNmM87gk/rM8j14ubvQPXS9nBGTV4
+Y4powa0MlLIK2REk29BvzLsIGVgiODZU1zp56pJNKR6IvpMj7keu8cSOJbx2fnQ
T4S28lHrife6tegYTkgQFDp126LckTKPqzuRJtIBTxJw/HdQK/2RzQ15EcSIyXMK
LaFeSpzHnOme69YQz4phcDTo1neM0Ep2OXaGgc7eSr+FQTv4np7BYujIpQ1W4kMO
VdmbdppLPeC0MZe4I92QUmy390WTH5kQ6pA4DB/ql9Ga6jQ/4g/ip3XPa807BHPJ
nKkSRIDOYlxxTMKT3qVrpqw3Q0y2Ygoobg5i+z9cZDRyAt/QG0AcmlkWhkhMqRB/
pnvsrts1hLyxJFNjboOpqQOmANwxfaneTuEdzQkbfJupGt9auwPHG93u28KFmZVi
V0msuKxs4dBY1TP0EpYmvhpk//EwnrEMekkyHp/gTMbS6HGbB4s2ZiuLkU2s15tT
NmdgqLdVdx4cHDM4B1aEuT0t1d5FYqWPeC0w6Mc/tAoFV7EHBuY3acKfy9aribGm
gyRhjdRXJbA1bPe0h/GVU0zVm2HWQ3DHtQDhcuxvAh4XjEhLbvuVUnwUY7Y5dz+e
L+DeYWlr3HS50NXHIDzZIOr2Okdkr/vIyaYp55/1AftYv2Mu/6FHUmO0Ke3TtcYh
JaS1Agk8CwVEme8aqT5Hwdcfyxk/qsjwVdeJIDpy761bHpExtGRw2r11Clb9pUBf
AEURIruFXk0blpFqnA1yc47FkDLrcgCOOv7U0zNPPHpmZqp0AecC0jZZF+9VM1c+
H8fE5TuVYb29TQ7tVj+ll7UmSrngwMr4pA3lq6Yl+4uuObzPtIrjHGt7a65u+Vuw
krKq53zvPzbZazmstRI3z1VmbMoxJsK9/nRR35nME9rf2DJoxUrNcr0TrquU5bIX
QkDeZQ8FCmNQRdfpylw+sPLMdAMi9vbmUbc884fSYCue6XFP38VMUAoOHCyP9SxC
r1W3THg4GISXKYNmGOXaRXdGImPZ2qQgHcLZFo1ZnLPx/u/uJAkU0cI3PYkQ9lje
mFBdymy2xqeZdk9lMn73km1ML8AJvaoQtZVRjNxY1sVmCZvBnWS+b8T+NkPsJKdo
bLT338iXHwAVUBvreicBZY1Eegs+1z/QdUI9Zq6DoreQtL/TqftugkU3kYnaVe5o
rYOmsgVWWrXmG4eDA6hD3el+IXEUKsLab7D0d440ItKwRaDidCylUsNWdwq3jCxf
TcbdyXZb2PCBslQ43k3g0Jn4YWtLIio5V0xiO9NBE0xMkjNMb5G8fWTvFiP2J0R5
dzV1RmRPoFJ1kXSN7zljd6WtJGcZEvIoHg7bbbdbV4nxqcCp5U7VnEiIW01HfM5F
03CQOgFCoqOFKHTGfR2/jauehwbq/fxzRMaQJg49eCyPBsFKo2m8FNArILu8rDhw
zPqMZZ1scC/OYgYHhtoCD3W64pBSLe5MM34dawQ8vbzitjBoLJGcfvy5w7FrcMpD
+R8beDwifuakoMebMc7e3x4PfgzdwAXWp0Gr/tSSgxF+Cp+JprlruAQlkVDjc9bi
MRBhJWVJNk6ohvQghvbHDO9yqWIhfKgtK+daE+0lwJcEGYPP9dJh1UBT/MUw8Bup
KuKeC6IZs4cs/IOUj/0QNSmrLcx6lvxHKlcQ++sdJFVPnUCI+zCV66cwxUUmeKH/
V9oDsVCpqLWiU1YEpRLjksMyUiBqLQwYkK3RVBNJm6klLzGwLacjucalJ1lreQoF
TFvYuEWXMVirSpzpiEkp4hhgL9xxw1Ji6eYfJIrE50pSxOHKF9vqoKXqjb4hwShx
06GpnkSlUYUigyFgCJdYYtrnSafLNv3HaVVCD3ipHZxLMu9D8xlwObs//lRCBotH
hJln3zPX4nQuAG4RRcDm1mW8ZBHCn1/QOvu6pSf8kWD91iAGQnEXmWVu6e0W7DnL
/5dyaRARJBn1MgscNUj+Lsud0Z4hQPVZkl83yxxfyjHAu8lZq7VHHXNAQG2pELif
fgw9P0PLB5j/T1Xbcj7H+JlE6Ht6ct4q6TUt1sszrWMAoDmfO7/Kbwp/T37MYuzf
lzMFgj/HSVFdC+PyGcuLllgQxCS26PLEttJ9tU8SRP66suDSuYgP39Epst1uoZ/F
dAn+jF4qeknwL0EE2KkV23eWdJXZahLCppvYSrwGR8C5ep0wRK+u/Y+0FTfqWCeg
Uc0pJTlhgESv5lEbV4DHawm9hxI8iX4v3y//pVyAQvRiM0e4DGIW5sOgtrF+ntp5
1Xx4aViP0ZUXeowbUutwZZTwrqvoz6OZR4RoIq4J0+R/ou67yy2hv2eINUv0hdnU
2UYfQ3fizsxOKCfABLl4whzTm8KPv5g3EWyo5IrWyk/6FIvMW3Yplx4Lp3d43/14
BYVnHnKPzh5INJA6jgj7LLygfINaT+W217YHOy+9zbyyw8pkfadka/ro6mT9x7qO
aRq5wuQXHfNTUvZbQBXEzgMM8/4IdbJ5AUsmNlIZYGgMzXqAsXCBFQ3qy9zHWxrh
fHy12/ElfN0jL+WedcGdAxOeBhYrUfHTdrdBnlEg3lfyQgMRyMFBO4MHMpop+HTs
ZxX5qILGl+gX4uw+BrQ320U57Q41tz0NxRzTPp8HwnyCvWnCQFVG3lJtay/5EjAe
WJuOz8MzIRpwzCgVybbLA6oeE5APeumRIESO0Q76v5FTb34ioMsnaZLeCPnUwi0q
TXLyjB180OgHLsuUI3ER1OwJTj1o0tm9le2zrA40mDNoRS+GgT06eXJS2+uIHQPE
9Ekz7BWLRzD2PeVziGSYRfojLC0yrDqXHHpIqOyo0MW86Om/hZdTxNkqE7c3T67u
PLdXVIt08s9nI/DV1BdElsYHBaV6evATfQnPAoJHcXdXxdqlSyHjEx/55ifv2eob
JDHIUUVe15a3+BEAEeqR+aj8XEVI+gGwUDyltjAq4k4GOUwRKbZetYyHWwC9Jx88
YQ+CXecVxPtd/c1TK45NqRX8n2M1DVsAOPg5Pe4bfGpMlz7sT/MibjXrjR5vs3bL
2JU6mQhD2Q/wW88Ko08iLiXfK3l6xF2ER3P1RP+W4945JhNAnAjDq9Va2V60MPne
GD03yHEK5p63u2bzGvztMu06/XGsjm4/VZ3eu8iaaxEZuKDdTD3AycUbsdQmAIgs
9l/ZWMSlZ7SesLHAyJyN+D1uPynwA/4/nx7n+n7hmyq5KVEheh3y960pVkSQhkCr
hB7n1olBWHZtVTiAuFicbpRY0XHaLbSFx6E8UpyYfan/5IVSqo0UHU7RuX0D1XBr
5c1GQuCL0c4YzZad1yZkP6f+iXxh1WZWNw4W1e2Q5FAGwQF0Mw/REtCi32tyj1Cl
PJPjfTPL7sZyVE722JSNHzAOXeTGyXeTWRj7+ywpzFh+AiD37t3E1xKnV+e6kklA
ASVe/kfDAMkp/WGmcuv5bdcATuZ+PGeM2pe9EJnaEnaSRVO4iblsLYR2y1nMrEXl
n/gQPvDLnGKhOEMKtPbmDfUB2UL3DQMRM9kDBKg2M7tFpkYd3xZqrUr3xSAnfUN+
QUB35vxbu0usOhFf389oB4uXtxChFkj9BEZD77DubrgxmIq4aBGevZwOgA2p3+I2
a64lUa/Ljy5XmLJkLEZp3jU3LF2tlH82kcsnMNiwGI2YVmn9uj96unqj0f7OQs8Z
7PTXGjPrR8XhdnmLO5kHyzxuv7aPcRjHLh9i1LHJ1eF4PN+8uZkm4T2YLIpxoCbO
yzoaM01qwtYg4pDAp08DqjNV06IeZhNmBxJ+zHxp78J/hZO0k2qwIqyyShvjtUq9
cdBsu6/3qtHSCRcZe/82CNut7CtpxydRaMoVoIcjoInYFp4jW6oyVVZclMK6gNRU
kVf44kDBsTiNBfPfA4bPUOnn2RCTsnu+GydB3y213LtNizKFAnsGhKBAn1t8dyo4
OD7MVmE4JAOL5roqhbd3VvWBD/YPdOLs3HTw2dDJZ6ZS+joccIUqRnX8ZsAfkPUz
A7Pu/vzyvk2yWX0cehWGCKuth47YJ9VWqiOoWYUBIMhQV8je2pZ3Rm1gdcaZnPI/
hRXSxlL7QrHEa8u1PiA7wqg8BNt5hA4vgQV1URb1EphRI/hEDWYGbPHQAMVC/i5a
wM8Cy5VdxFfG422vooSoYwXB4zB92l1Z7xYauGQCLVFj/Fp5J2bFWXrTJLvuEC3i
FywGfLHulBTwzF4emuSDXoDlCrRaj6/4EGCAmsEvuRxQ/Jqz/oCXwPiVIgZqpXTn
6CX967S08G0cfYD5F8nRim2NoM4cE1RuYVYP8bdw91PkU3V3JF5wHYa0MwIAXbZa
MsnMHp50LoYGYYILCuzKShT8oXD8noIk6p3UyhBylJVo9vXq/Uav55s1hTySizW3
s4DRaY5WkAFj65mK3gIFLeIpS4r/p6zPMre7BhsB212AiKuTBYdMneAGtSPmcKE7
OzeBmT+slCLOipJsS/nOUUYbxs3IzEFK6Jc0Z7bfbCI7vpiyrJdMPgB2dyxOqgGF
xQ6yyIyN5yqnRKnfVJLMznnxNd8pAlPgXyVvj8gpEN0LY6yxOvq9n+MjbN8Ayl+7
wRNOccabL0B/9ydFtXexNXVFuMM3n/inin95YdaAARaLe4QKFZeqkdqHYLhtJRVU
7llHY/J+4ADGNHQFkbrbrMwBBmj2nkvxuaTZPvhhRXEf5EiGRBHlTOiX+t32lP6g
frjpckYfOY+nGpn7tZhtXUCjXiAVkVUgDrSlOCS8hliaeke+mwTQ1yeHqeMXM6Dn
mQSMNrRiOYMGx3P/itBm+dIjZRdZMO++Mu6zrP8R72CPTB9pXTNrEMeyA7as4bA4
LBTw3ZODSSsJDxwdTWALCZyRlcK8zigzR0qvu6+ulkt4+WbzEHO0QjC9TRwJhoQt
SPItrL7JsO5bffayOOFm9JyqQ1Xq127GTYvlW6r4wk3oW5RymWH2C5ARssXtONTI
1ID9vvgs/0jItcjJ9fmzv/AM84ejSuDXy73Wfh02bRV3EWYmP+OA3ob6FSlE4x6u
PA/WRhCJ1XWiVx1LOrxVyk9kO572ZS6dDfkMyUafPd7tz0ofz4JfNOH9iIvt6RFa
bNJaoSM0e5iIeu08PpXWbcUZTZnnrl8yMlfJwlOTL3nzBFaoBORNgZgyNY6nMzIi
JyOzjhLsRE8vHq+QHrD+c81DqqiABE80HfovNi7gI2ejkHkRs12NrdVhZyXwopva
kOtvjMkYJVWlJOiodmHRhjkcehr7ZKt7pymxEPbmvOafbK/cKxPYCL7xLJVbHhb1
GcPliWO+5gmqKFnNXTB/HzzBDctOXULfp1a1YZxsRKnZy0WzEGlCx9MyGOmJcTu/
Srh4g/GD8lbPeV4wL4QhJFlOCesU39a/+OSRQKXRPGbtYHEiyb63I3AClhMtISmt
Lumq6bErI8wN7YjCB486HFrsjrzoMTa46AuQnrPO8/YEU1tCoGWeTeaOs8lPGVwL
re/GyNukmjyPtAwPxMpK5bPn2kTvSu50c2xtWT5Y/5P8ad5MTcjH1CiLrDbZE6Dr
e/6DE2B3yeomTE5BZ4GPYNB4JCP7KX0BJyBSdtsEFLHRR0QJcTx5XMzj3DKMiOPN
QH9o5ssdx50Y9a5qm/29WW+amqafrYSwl+SlsAk9VJMLWcagUwoC0W338zF6Yw06
xkHfEXQAOpdGVc4kntVpw+/7SZtvROOBRBH+nsVXRzY7Pw/URtO8CsPB+RTepNJd
JWw+7lFxUzlrxoEpEYlZAU1ONoeW1g3tGvuTTv5HLR9OkJ7m0bssxGYb4SSDaBN7
X+Bx3NMCPc/A+H4GVs35dR6r/r2jAQIMn0bsr7BRkUdZaBwX9g3J4s40HtdZXa1c
K2NmUmug+DVVHp45sEHyLrKCAHNDMcJLJU3kGXHiLNroAy7k2uLgZFpd67Dy8T0x
hCzQo9jX3iIbpaO49z2Cv/0tS8DW8difM0YELGnVoZWfLg6VRVxkWPzD9PX01wHi
H67iO+aeyUJZ4Eb5UUNXCbnq383Bka2aRXXN/nvXnWeiVHMNJRb1iFhIo/Yhx+3a
ZzA4rX4HZ2MhUIukSNDOHHHeEE3MjzlfnsEnvPNSB/nBZ2KbNZ7LJbkz5wJRuJhg
WzlNNKVuMVo7DEZ1vE7gOk6qt63Id54xgGs9bIS7lkfqA5CXddy+nvNSva++BnGs
vAB+WQhMbJbl4LKPMMsjNZUoz0jWe/jSqW+mSg9ngyW0pgUteoQ7GF+aX/IdAN3p
P7ogZmJoHVcrCuM3Zrns9AW1Ah74ePVoS9SvxE0517B2nn5UsTkBbIJLkpu8buEz
DyF0r4F0yND9kQxJf1hxqdtAZDkh0FaMXr53ssprk2LTe3FivOmkMXjpK/2sIMIj
DRUH9mCpEzydA0Rpo5CtUKdOemIzEwxPKSMyw6Ww8CMO9BCHtI3Rsomb9Jjy4q+3
AcXGpcdnAu6S264//XFP6hRHfP8zh/DZSuv8diC10uxykVRmo1H30o6CwyQ0lo+1
No2WmcOVrBf2QJ2lCL5BAbAFVNVU2Enh8Qe8jViX5mCGJvCG8gDUmdWZHCiOxIZG
xEniUpAB7Otvbe/puMB5DqmecMwOYxxh4qnnT3FBbSwvN1mzSWV8AwhAEnptmH87
39/EjZTOvz1dKixBmp2ZDgOEo0tQW9bTspM4hjuUTGchBbtaDvhogke2V/bOnyjF
QsNCzUGUDrntYlQ7s1RVb059p8o54oanXxA9mn9Kh+fVu+qjLwtn9E8gz5Pk6wzv
cImSQNchq8uTwHmRdjx66R1gRFo2dqL9S0uww83pRPDz6YBDJKiiYdIBC64klBCX
e2GVPcdJhbmlVc3x9IK5H6FbOrSIJAKY+NTmyLql+OWZgtufLFqwatCqSmiTqh4c
VBZqYhdbpjLwhG0nd0zguc8LVSFsvonKU6RSFG6ikUg0ypmVs8+U5D4PxkapNHef
2+jCJrppRvCdBOaLWGumKOY1WJZVIWjncuFia2Ytu5+/AmKzvADKZo6OBJCmDLMA
tMIfENzom7KbhhmPIdeiK2lypdt55mWchZZ1XPEZY8HDCBYRgfGNSd8c3adXlFyN
k4wU4QUjNkF2ICt3ABPW/VY9D/DGACmIT4pDD90lw/SVTk/VPjguX662jlESOJqT
xQS6jHBnDRBOzLwAnbheIZ+510MzWaytV3N9wVQKd7GlWhpIX1aXbFEgOT3HDcyU
cNziNeJHks2Ka71xe5/nmO4dZ7JOoPZJrSyvStLQY/9iudYQFzy11Xaf9+YMeLTB
ETdhkg2bwDx/jkDJi3iI5E0FAAddXFi3aDJWH072RWBndVIEycSQrBOu1T0r/Jdc
2NBZrhxrY3GhENwNTdXYSLHMGL0wbTGWwfJ1hboy2Y3VGvnIPqjI1TG00FtAzlty
Uk++CWuKz+qCsRZCl1nFUn1utWk4bOLh+eFFgu0ppo25Bn1PWUbfI83q453ds3tr
ljM73rhP+qrpqxcSdSntuHkEP249gryzQFLjXZaDbcufUh6ka0dqL0qjHmqJnLYt
B79EXoB32pwhdp9DQ/I6138XHAvX15eO7rB0I747wo5Uh7dtxyIVUUBi+JoSFXeq
yngLxwTL0LTrMamJ0ltPP96RhlUwSkLAnmrs8odhi1xGLMLo1WZUpzOCqWwIY3Og
yjH4iY2mMC6/gt3dMGEndLagg7zFzY06wuLfR0fl5CNoNy/Vyq3XDwCswmhLOpur
Zrf1tJjKq0zy+yfyeC61KCqhUzwo4hGYwnmrLnSz5SPKgiTiH5JZ1/7CSWX718mv
M/fa6jyFkzkcjQVtGSOfpSneepvGTM6t6jKqf6al5eE0Qtthg/vYWLhDuKEBzGtM
mBTV3/BPmjJeWDniQ77uQpr3wvwgsKQIvv+uBgV5v+od2xhvS5E5clrOMRDfOpwy
jgSIfrPZjGRy+SHdIpsNjR8g/F4pOW41+PHM9277uBknzRdt0r/Z1QABqwJ/etwv
ADZxZ/kJW8u5Hf9LglZ8y7TBjuqGhitBH2hVSAN5uH+R31dKaxVLD+hg3BPV7xCA
jppRzOa0eXnn8FJ5Sc60eDJ8ksgt2HZ+8xWQjzNidfNyvCxaz2NvuTqaLXKvmNKh
2I8Cew8yOuqP6M98w1aagbV5DqQccukgbxAqdmk1KwHLie6ct9r3HKEzUeW/k314
KZ1MBh8Bc2ZlcWGe8Y7jltU5I2aWz6wGcyYoVylMUyDG6rIE3cszaEptKFoUjex/
E0oboyFlXw98TvQI7WhZUYGM/jweTO6KditcXRasJUKJgWr4Wpc//mIfHbGmVcHo
6xffGAoPEuzzWKWWde2y07IxVXuY2wywk7BRR/vUk6PxACXJZN/8CsWgHsEtPRL3
Qzh1FkQ7DoRxhP8qPPQuRG8ouP4AMFsuUJ80GGE6rIEtd/ayXL1esVrTVULaSQzz
qvh9z3mASdom/D38Wu84Y8HWEDvC610eQt80Z0E2ALRr7knLO7PJtrLTO03WZgNs
lIAFRRtpu0+UhgzALyRG5D6JEOSGLnmU7rj0v1G8D6kkRmcbG8kW3EsG8jj1Ze1v
jGOwIc9x2Ljf3fEzS4DG5JSnjaM/a2ZwEh2Jwlkz44Aofov6tE+kpZ+HyYjDa7OH
1EHiiVC2datB0IzRuylSwYCpWEJOgDHlIrvbcfULcjAStS/yI647gxVq4k2YOqt4
lg17g7X+DLqa+keAcd1qkL/1PTh9Nc9SR57JMqa9a0hydL8mGT15SZRuBl9j2pfl
JZ0BryoK6AIAODTUztym18DeT+eXjAcfBc5aqYvGLyFzvnhd1igamS0OEfzhABz+
OLCGHkdkcUWJJrzzVQQs0+BFT0stHwygwa+hATMtZv5vZtrLZ+4GNRE4H+sqauJl
/m8cSPuxZLU2Ax8KJG2A3wJ4+DitNS4AYViYecyDzj9Tdvkym+NekfY4S5n7yDOk
CPRFoe2EcEeeNr76c3kg6Gy45VXz5ZxDp1KEsnf/y3p54zkrGoCqL9izKN1V/cNj
+qVUg3Lh7gvWovXZarrvGmmf6noOaGRwVCfh1jdnK556kYdVIc3J3A/BEmwK/Aar
Q7+efG/twCONUA7/oi8w++v0O1HsxoW4VU2FYDS7NdNkWmAYAS9P2F/8czMU3ckN
3fWFgl1QARATTM1/Pxl4fl5Ri5Etpuf5O2OMz5H5lAqieh5Yc8nLm0OSMI/3XEAF
WqfxUcD+L1pa/qeHuNhJZiUKWYVwOGTtmyBOjtfg9cFYQiw5hbNfsbdunXHnCCji
dHDtXCVLfppHP06OGgfCoVaCh5Gu/t11BDytOp+rkJer1kmWQxp8bpPM1NGHwr0v
DUEvDDB5OkEwlrITLed2JTRfoVXmMozdaryujZIw4+Zovn/wmuJ8dvtAiKFqjkT+
vdkyQNm2JjLyXk9U8RMYqp5e9+uyGd6sL+oPw6FIyBbSgr8pMgG3gzx7NYy4bEUM
8vz2Q2U5JKwJ19s1EFEvLzuhdzxnTx6rXs5Y21pE9LI460czmly6yECSK329HDmO
aOjp4YpeYyhjFj9G/FpO9d8kzZmMxL6vdxmD7lC3d1bLO+T5RZ26RRudbsl/EbfN
Kt+ku7c+xncKqcPkyEzfnq67gD3LKYTA1vf01LYDarRC2tHodRJx9brsWI0sR/Ic
letvaqD9cn+ho1CbUmItBwEh6EwH3VY3RFEMkWHxvkmAeClno72KVCWf95R1KkMM
YRx7rwEeVE4Z2ppz7COZ/K7dqFejr8KvNxa9q5uDIbvSTxhwTsXIMLXuntPpc1pR
wUrPxQHE62VC335TpJ5QwViDFvch6R/oaAO8S4BXHhrpUlbZjhFXkgGXMJkZM7Tx
8/MeCw6q/9Du+SlHyrMg0Ks/sFgXqFvSg4BQG97py5qdiKO+rWV+NAlERApfP3wz
44FudP2nP0dvpR0NO0Asffe8fHdc1pk2ITSnK9I0T3gBeug5RYcqKBxPzhKnOAXX
vMgXWatcNjF0Yjg588D5rmV7PVEBO/WojqMxcLgbjV2UlT6V8G0CJ0smdOe4QL5/
fBbPAdOECWjNNguujXB9M6kBTMIO/qc3P5Ptx5l7noNiZTX6lfsHpMW2iFrt9wvT
+BotRM4CCVSMiXPeT2QsSaYLrwiREHpeKTCrq56m6Vo3QTrqwR1snoivFwMe4ftP
IFx1DDnXla/KjSOJs3XO00GVxT8KPI473CxdRazoBvqVe5agp2hsITXsQSHD+MPs
3ESXnZ2dXKOLxRNC9D3Yx3tpYvGmoBtt47BgSqn6BRrOGUjtA2rO/vFY40oku8Pa
BDeKM9bxo6cTfgJPZttH3ORShscxdTUa1mbyBEgZ2bOvq6MD8iVtsPfV5V/ZWH0v
UsvrAY3wZ92tJm2f5iKCfotsupiv/haLYhIvswZlFHo2alN45v2VV+8QFvaVjobs
/PkpQAe4G0+p9zq21YAjgkieXe/ZOXVhzNocJIzDYtG1UDEt+XTL3MNeUSFCyipJ
RlqU522bt1UWvLutJNJZKehSbdExnuhh1J4LpNFPAtnaTsTWAuaCpZL9HEtAM7f5
Jtwll+/jSU2PuLCcKKKJpHj4F9DdMQ2isTbb4aKzPvf2Qwo0+zFv7ncJ1pTX5zHd
CSI+oMYDrHjpZaVfsM+/HE4fOTd8itc3wmewPY0DNR6jSgWsjQNLV6j63HD23aBL
DuxXUS8+TrI+rXD0ndvT6xAzJJKCFJc/VwA3LkEldL+CWhIgQZa0SfxsBDusYMMF
Aiw8PIdyLYBIdquna8F9R4FDtJvRc5WaE8cY86gMSoaZsF5mj2DaeQImjYotZgy2
NzB4FPhoRocc9knfo2SCbzsE2bZ9dq5xglawBRmU5TV9z1DsXMBK1JaFyKT57ukr
NTjiMEbrOmaz+VoiL+Q0+OamIP0vhSAHZLWYpeO5XX4uqWv27AlEke6pjuS7tv58
P7epVfBfKzSls4400IBUdAjvwhz9ApbMkMwS92U3srQHGQbSDAdUSFHXgJ2bJF1C
afJE68CSC0NvIpo+Tdjm8DBCToH7nLjweLVCbSaZsqYSEj0wcPU3nEfHJQo/oRPy
eBlQtnsq0VP/9Mwm9cJgd1Ok+IX7IfmuUzLaBZFFv0nd3WAyK2FI3nKwwdyoCLFL
MvmOAw7PzyHp4Iw+9RaPwOKucM3Arw0pPygZeMsU2dKGTcqX5VRsl97CoEjsuYcs
i37mwLcRemWARSlU3npdWPegjmy6iXBoNqyDbMpTlIjmdCnRlxNWIwEu7hAJdqop
dwtNI3OqC6OSRQ+Ayw+Q85YWUzkQmvp767y/DnGk5FgPdgD50moh7IrizuiCMn73
GZL2Q7Qcl5jg7PQl5aZWzPH9Mo44xoAb/ICNi5zvFTCoEWwLeNFs6ymCY4ob5vnH
R8H0HFnw/2CxNAflvy33ZQaGwJiovXm8rPkRyFDDNXRGFcMwTOtdNygktWZBMCo3
4hPh9zsW23gHlA5CRt0kGqBwxpynwQTMOMbdPivgq6nJ9ibSXS6UjC9CU4gm6WcC
Jl/3f6M74hyRHoLS8OkcZITLkMDTnn9WVG2gkYwrzmDIt3622Jh3E9dUXK0YPf6w
7rb8+SCFDCdaYWhJR28zdZ718AGfJXDJYv1zwd5dsCW4UiMqpTwEf8Ej6mObT7Nx
2AUB7RIOIhbkOtiyVjn7kFH1XUhb7H4FfHhC6YCDPcu0PQ927JxQwPODVxUQ8RcU
1/p+u9OtKRuMzbwhsREaCba12mwiCBrDCjh9HREVdZE6YB+mdGJzvoouSqu8D+LK
GxRiKQ8vEj8WPOj3e2cFRK7grYy/gXVROhoco28YDbVDjNjy8LGiYd1zNnspnva6
IOIAqGXbjWtkntYSpLz+AW1rP26K2NtzKbee8xJqkE1HfCFX+Ped+Wisn8P6uz3j
OeOc8l3LzqJ+wBPi1fZKvYF6qSR6hYSrjEog57rYpWq3WLWtdzteFVZdnajml9yz
P+XhnABXjgzhZsWW81KNHi/HN+G47BSqP/hKh4tT9mCk6b+vETHI5JDBB845tRhL
yCM7xHiYJcqw8NYTKXZwIRlKA1cQ7ZxC7+TB189YzXFIAzLfhS1IcZvTqchY6S1I
d+csIzH4demxcYf8Djkm8mEddHUjI6LnKI42asbS2EXSAsZDC8BsJbogwKwa71Jj
hfOlQw2n3PaaqzhKXSPSGyie9NDOhTqjMaqLJuKjODTKU3iIF5jKWAl0liA0apcT
8mSMNeGTSYOWtUmWUyGm8lAMFfugPA0wmfXOIG+8jxCi502EGGqsGLUJz8Dg7pe6
bqbO0fbWLn+Z6nPMbVJ0eLxdyT6Y3oIoIjAbRB0tgL9ov5VyTzOtvPlyY5l5R1Id
MjYVu6is2CPvcPQayvt77semyJz/cY8A4xMJVzir907FlYs5gOYsPzXBII3u0Apm
k7tvlE7qaKw0/1DakPZL9gc4biEtdXkY6U6zS0M6e/LvapIkrJU1hKIi45jq0lQ9
UdY/l83iNt7qdf4u6vip0t9vkdpw83smUXq+jf1GLZ2wBEHApCg7K5e+dx6J8IJm
RsQ1tNt3wb/sXiWW5aXCtQh8I7Lyp9wA1cf7tXdzuMb1htLxI9cDjyIdQhJ53Yxo
yAsCAOEIh9sMQAc7EUQEjW8VfjUItqe161MaYDaNwUPhYPw6vObiNe2UJNx0dWmX
xXBUQDiRXUaS+FsqgiCAClr4Rp3DXFfURwxpkcnIdF7lS+DBp8QkRFOJAdu9ZDmR
PB917a8rMBbMuzjL4JgkG12oCUGBLPfmeqYVjIUPHebiTdQgPOnbUZitn2uuVVOw
3LNznHlB0yyOrjnsHaK7sgyRV231r4SoONWjVpoM/rQpFCgrcPUSXHKKsnGaaQd4
cWCNlM5mBXx+uYhv/5vqaI1iFLKaUFg+Zb8EiasEVMWxHjjrR3mEnPR9zVHuki6y
Nw99rHoFFc8pQ9TypcpEo/btTCpCk02gPaLbMCAkn1vwe334A5f4QPT/8ta2B2tl
PGOAXEvwrS+hBog7/JGaGSJmtujlUoKI+7bbn9JXNPL1/Qsql2sfN4iwhnxc/3w9
eJ4wL2/iHHAyL8EGm0Ur+EkQ1wS8iJJnGtD8TFi4E35Ycfkrs8BAuudKPUGQQyPR
0mZfaGKbm7elwza5eEfCzdaV3SsgUb7F1Do5eER4KSn1w50Yvo72MKQdybGFd30F
/5rvL+fGy7DqYi9FJqFtGW/wGUnjHrF8YqdmEI/zgDnwE3bO2dusAfDdiY+T69qq
14GtEuRuWx8laAa0mJsBnJdCrGpvsHfXRVPFhQW8vse52hYBFPbJcSh4xoGaoNqx
etySBhJtUoYqBJy1RxjermFEpzy9MlColWYKxmRdbYnJHMLbpbUm/OM5ldH74I9T
9pnv8/VX9Hw6Wo/RhLr/WoXac74HW6K6cBDmXtoliYJWRWeuTzWzXXah2FhEbqWa
jzQ7KwDXt5NGIip2eBoLgFgde47yzbItR2/hlD5VW1CYeLTvR4IgbvIYk5s3kzJ2
gy4S9SciGMSXZuPYAVgkR/3y5DjqCsW2Ru/1eUrl8qdKXQwU6xD+IiI/GATyDFIC
FakT1zw2211I688nbCwFK1B9oDtNc5rPOh7W/dI/LdKyRDEWPntSnsfStrTxlibJ
oUgPDyqO0uXT8Bo9LZiPTt9PnXryOPqM2LZDrfhpAspEOA43pjjoto06lD7S3U80
ttYiXwvbfC7NMCxoIaHkUevBoWysNaZYoPECyAJihAMzByQyopIdKA2iTnaMsJrW
YRcz2YeOqGike+ThY8elLiEtwNFNr/RR6njwOc+qkt7WM8WH23r/K3AE6mv/W50S
jKK0n0T3vxeI1po3Ikr0bJ8JeF5zj6i1a10OfAJY88u+LwKjxV+RP5qTQTCDfeZ2
NxocOQ4KN+14xsnR+2nbMyQNMjwPjjFxLAqXxhU+DYCa9xx5YAOjVVmNlvgB8rgq
psjqaSrCJAvJpydXij7hNXco/ubRc8m8SqfcHF3vAm/Ypqs5MMOwPe5hdJL4u1vI
7BDFqBZA9JFmYs9o3lb0syzN56BBYd8k5uir8nVBxfw5zwA63yIngXI0+YalSIvL
EikOZIQ6V5BL13ooqds24GdhU2Y4/PUoBjaeHxeY5Aod31cYuqCzxrEkgIHbNr1B
ALvtXwnlVp+S5sFsisOmGbmDZEkDdJjJjLeugG7HjFPR6StYzXvswbJW7iYiI81E
T9oTtdThoL0LFW+dmXsPbSi5ZSNSMB7trtGCBVaR3Tz0noTGWwZKktmomAnK7UDU
pKc2ceGzcFoCF5zMXo0TjB0K3RkG6+WGyfFAXBA9B64+leZEMlve8eCv3jUKPNuQ
df858Y+54OPea7AqjvxTh6EgVYr87nKoE1BNKHif5C0nvmUhq6ha6nMWiRX9jkc4
G7/XFErA/QbYg9PeRqiOvaPxQyZiDFI9IbvrIkbUg9O9NKbXG+UD8KMw2s1L3DGm
SiS8uKLDIPFgLUXaCQ7Zd9Nz6TUCzb4BJ9gvTykOdpyQVjT3d4M2hV9l4kgBkcP2
HF5o1sjpGR0aXxBR37uQB5MbQ2n0ILRtPcwsebPZMXg1Ytgv5/Cya6j6jhLFjERg
yRCfRYP7b0h+DJhVfccKYUDAj39brdvr4cA0TNngNmvaQQoUOz62m+Rf5k9IgWsh
1hRc6W+OOLK+BxBCr7JxvSyJapxOvMRGfl5mKMnqylo5c5NkhIi6q/VZ0rvYKfVw
gAeEm6CtFN5gWr0X52r8Oj17SMko9EW1XJz8tVD0PVX3YdKz3gJ+aWKm/JkD1Ydk
oDsMCAc/h3cgEK4gcE45iBd7hf/7i8uFQwugVss796tu5mt7PQHIe/47hiEswUhs
BDEgaMWQHWp6bNfpcEW7WBNYDs439aUD25hS5bGa/LiD+6n90UoZXekWzJnN38Dh
qDa+6PR4zuXED7ky+kD/m88pDCxymmigFd0Mvo42nf5kAK7vfRgCCYOsrjQK5UtX
v72We/4GCzIay4tVn1vccwsph7rJ/QHNQCd99de63dR8DDnmRxAo5Wp57JyqDA5l
HtH+f45kbz7h9FV1NYolf0mdyOGhhV4HSM+FwpCs0IWIOomWtn6cp4XFFDbV4VzR
mouqHv/0zGr3YG+bYSYMRWC3SPcN59VcgSyca/+5VIvPKBTmS9oZoFJymddOH79D
eOOqzynVmy/kWMp4OzMv8sGPMC3auHwMWMCk6P7Rhl/Jn2TkbTGFToDCeHo7OcVm
+tGL96w2Ck+qYAG1X6w54bYFXImTJWIdX4c8/OpgX+gHzMff5GHmxR+7YY741PAK
XQH83t9U5JmOO3P5s1ZhoAN4AlKN1E38vEUjT/VHCk3aCAtvfYRW6yCqz8jdIY62
eLOgYTqO76VysfbXQu2mjPJcNa+QS270TrNF0p8DlysQqQBs3Dk/6RU8mw+YVLHI
2vH66mQR7r8VmXCa5bOpkg0f1ONBFcLIJ3DoF68e6GXSRmkoTX95PMGHAY1XpZ1p
dGNGhY1DPtLr5AAeAtZ4l3QToWIyxxHm5LcAuxS+Y6wiGyXIIj9Z6UFO6rP1c1Gz
eTw12X19Eq8nmagz/x/y3Jlov2ZXNoToqy0kBvaNqTO/UE5aOGVm6EFGsD460A7j
FnmHW06t3/DA9hCXX2lBri8wqpT+kM7iEBlxnZZDpqjd3EWNJsWMbX79pIwe4nmb
cSuf5ANQ27Y++yj6WsB/uXh17HkZ83e2q02a3e4Cvl7oxXnrhXxd25Xt4qP0e+n1
RtQFxWAsXU7MOaSv4tPGnL7VHm82nOFlSYNkQpbnNk66PeKyWoICP7sj7W7/cO7P
+cVwHtUQO/2gJtdZky4opX9hvl1yRtb5aTPNFTXGmz1ZJB8AjM8E22V/sAO0V32L
FnZp2JCtPhJaoLeYh9/GqnG3DAsNYv4mstn4HXysklKXDPIQut7BHKLEC6GfvdKc
NS3mKzFKWzUeGM9g+qJXNKSYficbwBmNsPt6Oyj3YFKk1trXQ344Uon6aIIiStjo
//UCysNw7KWfpc+RmBcSnLSpzoaeG3ZxhY+D96FbODSUKcg1AqcCgBucbjkXtmwH
JZHYVw0z+o4c/7ye2hTyAHMq5hYPdu9NR4ElFKbaKyMWdZMrePy2QOy2xn9lOZOw
fgHrE+Z76QKdi6Z4qMm7em5gVvQmTOAc1uB8Xkt/KYBJS0YeA/vnqoHfoeogJwtr
NIg0QeB7wgMaMBGzpcCWmd2cQ99VzocrNEMUN/m8Lsc0QnO4jGDeHWU2jIafS8MT
1PeV/A/W8nVxdpCVYcQx2bNujmuCd8Kmw3R76XL8Pk3hBo+bDt4fViZ5XY8Gaijw
PcXwQyUdJqM0/dkxl0nnLBg/QPcgxAu+NwNkDyVONSjKL47i8ojyXk1vESlnX6G1
XyHzFYUolgHk759Kp1fxBNgj62EmtjPjC73yc4OS9l97KQHUj01rfGimRnMYJoPn
fpOAy+Qdhwvk2x/HHgihjrDK1dh5A6WE1d3QRiIgoPrxM3OCwXd0LKdBQfTPYVlw
4ONexMYISNx9tN6FEjwDCcq6O3p5KGr+beWpDLIDL3xG3VmjkkiZQFrGFD68KOPH
RwIJ8HCJ3nF9BiVycGkBR9L6D+7mC4eBj22jphSUBnweqhEm+OO41yLFnJt8FdzZ
pZXZ2n2O3nGyqNRb/MiTlJAWgYrB+lfVnp8CpAbqIlVwjIxa51XO3309PjR1sTPE
DyOJRV3ApnIKQQQJrPF+co9SIxkxDCeTk655WQa8irJ9X/Or4Klj2f0C9EcPmNPV
1rsUZq6u2RDaoTklfpTUJxijxsc2XjVr2QBw/hnyC1uE799gxkgABGyOn+oq7o03
iEaXIuSc9OPjLFVp4YssKHxHRY/9RSdGZrZzJtogLOj9nbSYPoDeoXPCf8KJGRNH
e4yxYaHwgkayV1lQKFU2kc3IV01jEk75OXyWl7GqjS5q7ehIm8ZyJCvH/OFeSX0H
LNAMy/RzD7ySTJp50sfr0d5oJLDDOHuhGFmUc5f5VaFPhz2Rr574Y9Qr79qxsC4f
4P0RJm1hqg7b/7loVfd/6qzJajtoY/nvJfqBp9iJ/pLIvfuCCTrE31vBbjKEC7Q2
kPV8U/RpfIJn1/KLbHDUlw+536hjigXBX9m0bwYdxwtAU/cqgwLg19AORRvcDE6p
2xlhwVvVspGfmGMOg0Y1W4TNF4+EzV0bH9s1vOBk9MsyRTUcgq/5Tw/4ctjeWpeN
C9QykWjABCfYMWo/7svZLSgjDqZoO5rP4bZ9CIiB6BMHDMKdsTLVzsfhF2bgP77B
XitpKKHz/8BQT3TLlp4gvbEy33/C+Uv/pJzKkJ1DCTDzYZd248fYNnZpaF4zsXiB
zz3UGgAOoOaOAfIFzmNf5cpqQit92i2JAUMsk9FgRZCPK2/XHrqIz92FZ9fbO34C
drQnmTYZEKDZFGycvFdxGKZdf6u8I8pqY2t00Zj3GUQ27ffS8AoKegIB84GzSF15
ak9k2klCh1/V2TOfHLnBSrnzQjXyAgG20HA9ImNubEyT/5bhAdXIUJD6o93idIO/
8PzibTB69LUiHDmuZxHiHdD6yuaUn0IyAiSmCSC6AanltcF6uWyonr/WvV+n/Dcp
lJm87YsgM4Jl6Q7C0H8QJNB1CP29vDDOPKK1xlSDJTbqljulBCr/p/j/dwTUGqYd
GEnNV9tAUSKRSWly+La+LAV5F8Z4KE80aQ68H8mJZS+gppHKz9uzvxcTg7ls7p0m
3JIiXORxONfFw524Dz8ptwVW2QhkiiR1q1IcIHQE4mX70pIfkj6BAXJyHd9RGkRw
hIHqP+KvADgOgiWieiJqnSswvkvuEpWBNoGBMsNxskOBZhuOefJRZ6xOLnCGbFFK
wJy4UMXQUmWFklBzCzYRmS7P6V4hHhcnyC9LgwKMM+H262kgqVlUP2vqJx8IrcFK
6QrcnzkIDz6P79ZUC6pq9O+fN10BtRKZfOUlcDnRNJ8wQUtgQTQcO89ozp7u5n41
xuIdqZErz4RrVtUBfYfDDg1vyj3F0/4YJSvaR9nc5RXPljVWb/qRHsA4m/HE+EDf
YRY2JIbw1hjpv0Dk4FlN83bd9lvOrqSUsBUNvJba8UHrlrzSsy4RImdawvG1sl0A
WWcdBh8oGzpQ7AcaxuFroP0DbWzdnFzG8gAjH7aREBAbLcu5AAwRrFmSShX9OSNR
MtA5pcqKBzy4yurEfRXDXU/jaRaMZAlw0w4pbESCUWF0vZZAM52sLQCHB+TJFuim
OYlKws1+B7/pCW2BBii0JxuWAFhJ2TmDOnHf5vPdcmViwqP0jzkMPFayuBVNuEsw
Cj5vW6ieKg30sCls35qZ+whGmGTJyMBTArK6gJ1QZv87l3GdiCPOdnrAHDgonDAG
k1iNArk2T5cZRQw5QM0X9uHPU2h73M3RXlByIEkF6cmpO2dC8oNVv4p2afqIZzEf
qjk6xSp8ks0jORaq/uXDxLczHj7BxIBzoJ4YFJgtHGHo3UZ9FrQfnVfA7tkwGAeu
nw4sDX8ZbzFiBSMSlDGX/HBvhjon9kdUxt7fbgww+R5kWGI5FqcreE8/siWS2n93
6M3UEO3rSnaIMrCSp4/D0shOo+Oj1xYdYgLfMgB7LQjamNwQuh4jKFf4UdO+o3LF
p/iKMfdeg1Bn3XtB9NvuhcIp3XUhN4JNUoBLpkjX6efKycXrDiLTxH0oFZch6CaA
E4zS+ZrAM75nqS0qDbYMdsqkeOFCB8cefgFFniovv8lTy7un1sG+S2QTEaeWb1kJ
xi8tbzBIOyDi6N5nwd5w2NuB488Kj1zKeI41fFBZkfC040oEECddSA+PxaMlHly3
w5XGvsvhngPaA/SkVK0QSc/Kz0UKFEYGg37P2dK1PciiKdKqIQqrIf82e/+51Nme
7v3SV66IzbYmus6iPZskifo9B6G39FHgTULfckSnUCZQoRGaQxGk2U/g+jqcHg5c
tC7dbLQVU7CpUYuW3BGEdxCDoGhzSfvDPvAeAOK8NlcqhDqOaD6bvqbFKYQTndUn
YpDUzlBbOJqfeHKQqdyb1j/ssQXX1sLXzuI79HPQm+F11xRNKlbxTFcvhZgzu0wR
vc4b79QAKPTqQQ/xyMJR3N9n1MXf9jWQwkveevhrkZWSDTWfZNS7VDL4GjF8Odwi
CSsXQ4F/cgH2ZIv0pmdammiPigfiF2yFQ+WvOrf6ncb6aLwWyfpKbmunAaRCSAVj
9DwilvLAptley481+gjmrWSAgo6o5AXjLGFO6I7rfxY4yfIWermB/kMROMGIAcGS
dkeFRF2m2g6gBcFmLrGqw21tws2F9uvSBhCkQkC/vgDytrT7zUZ4P5JseddqUIRw
sKOiBDuM2GPE4rvqg6a6B9K8YKTog9+Ek+30tiogacDEGsgZw2lGHVcp3px131iM
joC2yx0Gze5pbEd1labUw6egoRC1DZfEGL28AcU+BbaKNV0HKW+vmnkGPKsjauJp
rlVh7yN5yrvzkEQClsWeS41mzLn9VD96XAXy+xqdGLgSyo8vL5umVMdJMzUTfLYC
Pvt/AXiMrruSyFyDR8HCORWQ/tGJBxGX2Eol2Ffgm7GpvK0435ii/pojdBk1NaS7
5m37f+sxqW5su1MR4Imp6TS6Jl4PdaIFsSisxxINrk88FbSoQtRyT7RD4VuwzIsH
+aY/hOetgwGRn0atWYh/+6WkxB//ZdGhmq0qE5rzpeBgzuascZUTQbo9zj+FsPHq
SCoIwGrwH4gMfg3u5BFv49Pry8Ncg4QYNXnuexD8F5H0/lsY3tUUTb/RjQXNkn24
psC69hJmHb/tfRfLMm40j6Yx6WxUfIErJC3bFIwD+cADHWsERMigMhuapDFzkaig
RUjx/GJ+0MFahfzliRvdZgVg1KDKicrZzu+fU9SAUDCyfTdSTWCsQx15u/6NuiJt
aGHUdWqS8oIN1vtzhbV5firj5elEE808Z+sRu7opgezzuutbvcB2nkn3glVS0Sug
sC1ruWSQdsmBFB9fnhhWD6qNqwCf7FzFqLgS2sKNDm5du92inNPlT5ksg6hEjYxS
AFv10empY+AykHI67LwqAPPyyTxPhKCFnzPWeOMSdNVX7xENwCDCPaqUEdTrG80V
oY0/DsFR9LCovELkb8VIiwmcqQFU/p9gJZP8+pEWLbAjvAjvheaIDXaBX19rfEAj
ZaeK/20TYRqVZQ3e1F9XbNz+3UHqRHKbGTdEb6KFtSvXp0OuGvQBuJpMlEABMsTv
VIfcWXIsEWwzVbyaTAojfdI4F6FZk1oTzg1iPfxVuaCYMmpveObsv3Kt8bPq6qn8
wVZWU0a5e2TXT/g/Gfiim96yA1LvrOVI0i0ASDzzIin6zpGd2pheEL6IjaR5yStQ
UBuSUYY8Wz0QuNHQUTxBqhU8IVEQdIAfRIWEH/1wikEM6mDtXXOs9VfjzH+vbMNQ
kkIxahE1ZFnlRBRd8hdZkwHWa9qNrEXKkjudz/amPJSRaexmJESOqfwYVqeaIW/e
9grDZFFwAPWW0MVXCjtPSOkhJjo+WgD7FQ7TyO5lcdV5sVdOcPvmTg7lihTZKSfp
c/ZFHQSmf/7ITgHvQ6nkRHwrSGC0yb98FMaqfDFrdI5g8+VaXCXeOdIcIrInpSmn
4PrAtgdUv65OpwShGXTtVQpqV7yEIBvgCPtVlTjL5sXEvEqrujRURJG0LDvi3+sU
4MkYKN0EZNYlpQkR8wyNbM0vsErGmgBVMzKHo6hVSvcRTi1y9aQsHpnCUig3MGJO
oKNkcQzoOjihbSH42X3l29lqrc8SSEDiM/dSBkCFic0QofiLIww2UU8RSNHrYfbh
FXvsMXErzUy/8bpB9+NJZE5CfrsvRqYRqUMSUvUdz4a8iTqjuyMN5znWC/AyrtKA
dhjF7o34B6Sd6sXSb9zbkSXiloKM2w/YpnpCe6oypUGMXrIL0WJlgmIdKiGsLnSC
q2SszWOMpdMAE3Y7SKcV6A8S+B/DLc4hwpJUbUIHiQL/bnmuDLdET3k8ef8bZXPf
xLjOApMhe8+hAZdvbmbpwoOmJBDDtiN+ROkyCMBK51IwNTo//yx/4gTzfJ40Tkdo
n9py34wgeT66KMq1qDJ5f/5WR7R6zPZ6ZfvSV+HKxAOwFnqshSjYyFtQgDPt6Sx7
aH998k3fmKnuK6wB5L0JgKmRYG1Pawn+3ks1RzOc3ohLcF5squBbDLEZF8ASERJs
fHD2HuuocI9jXYWzvyM0E2vWG/06oP4OysohQkgkKykU3ji5dq6mvpEbPMeSW5o6
+l+J/s2KQRicz53lME9pIewDtkJpgd2TJ2AcucKdDYtMumcBuRRJakjW9ewY7N0M
aCoFm6Doy5qj5EpGDnRGTIZ5En3YxgpjyuQ9C8Zg7jEBkJ4ozbhV7RBuE6S5XNIJ
eXNKejlyCMHHAm2TFlHS02311VmptkE86ps6myODicD9zz+Czu2Dd1KPPlc1Lk8/
7jhAQsHQ0xyWk0keObEz5RwAPy1DyTekac535uQYasN9cGyyM/4NJx6G/lXEw6SM
VDLmqrU+jTVhsHZa/DdHYmQUA3XiHGfHgbQt/6GylDpKFE8KImSpLIIixcvSfYIc
c4WtXnLm6+fRRk0c/gzj1+r/orZi3zGpyCmr6QWXrMAVzLJHWMOReOH7TbKhbe+U
5M5z9JwTUmdfrcu8CsuEXb77K8FBVPrQkkP96jUDqZp9Rk1rfMWbG4Yv203VPtb2
bxtv54EFmNVylgjj942VgpjVN9a3dhfMOgw0MDwXwcLUD6rbbFuLzJkt2XaElNZo
GOJw/B69nMfsUVVhwb5gGjfwZZgsaWDMp8HGm7i5p6GI1+kEMumQRLXRm29tPrm7
iVHTgxocqT6hrUjkS9vG9B/J7JmwtNDbACMH7CoWjX3zJZmO1NlD99zWioJy5BRQ
KDY9W8W6yhfb+AurY25VKOLefw14bpJg9893uD9iLbHeZKfmVfHoah9v0VEc3k6q
QSjT4dI8SuAgeCmzOlrzG79mWk+vdq8vK/cknU4CwpySWXSxjn6XvWcDbddR7weR
bQiC0k6ZCNxF6dGR3j03zvB8YEnliH80UnOnHoPeWbYYORkzGxsqNoLT4lXOZyeQ
9gyk7Asu1mY2gW63O/IJEwd4KLe6WABFBPCTsoR+DAZko9+4USMdHAYyj9wrZV09
0DV76wDVzkH08YRMNeKfl0ZTsQV1nlCsVaPZNfy3UHFERPN5+2wnn93VNHuJ+YIZ
z9107yxwwX9jk0gKgTLvyPtnq5Iyfi28RZCMZ79bOxz0qzp4tZkoMQHYqZEF0bKR
bOVSfhNyesSGTCQdCl/vlbti5bHvWZVMB3wlRs+zFYQk1AQ0IA1JHF12mbbahPoA
moCQiZh0b7yjyDdrBOzGX5bezadZey13ALhBGQp02IMhUgYAMGoIi/GPynHwXhMP
YrmRGycc6mvhkmsh3wTwaqDL7A8ORZG54gix28nTiCfTYjkMzCzDdM4TAks0bwmt
PReE2qmH2VgFduz9NTPwDlfK0tL0/g6RD6RvlFmIolKOeoVrjOshcjQLqXj4q+76
Ah6yRnT7/WxKXGyDrPjmuqr2DgWlc7S6LUxpXE9Foq9CaBheU+7dQUuayyeXdI9/
AlylmDX6KUjTbheUVe9mqUK8Wx0hcvd7XF/cmhp9HG+NoWPnRKMcJTldDRpYrQo5
lWD652c8plhyA3fW6RV7iQ==
`pragma protect end_protected
