// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
sI7aSw58h7UK/wmm1oegXrBNGG8tFCbI9cGwuUbclyKtVBdR3EFwzmWsNS1DV+q3zJCfz2o4HgwM
NNrOGZWOKO664f0hfIUOHoAXchlV9gJMuZ1RmBnzqoEcgtZuzTfaUEmsOMQDLTZSNUIsmagaChcq
RENx8aJK1x9rDEdrWVghHnRN/qM7iNzebp8yXhf2UP9nLuS610ktctXXMB3t2n6InGa9gTHi6Wo6
j5oKVv6t0xxCag9ZER46eO95eXMji3V9Uf9/Uamhg814lhYa6jyRHR+IQlouYmIG/w7WzRkLvPtB
TqwoH/5c/KkLAM7jFghQ9HVMot5qXOzv2FrqiA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5488)
bm26KR3dsw2hz2FWR1Uiit/p+gfbVEEshejUig/+qqyV+CA3MXAL1WMHiPFE2Q6Lk/AaE0ceWpzL
TWavB2daTlUTzeVxoCZ21NZdEHYg0F93eMhcHB0PfzAc1SnmeayWtSsfttYSQWgdq+PhFJN4oWyO
oBKw4y53HbgCISXZgmV4bkkWIjOzLcrE7QxJ/VpdG156BWNHJCRpo6N8/YsdHTOoFD7Ydcw4tFEz
DhBsNioxtOlrrmSNM5aDnOM5p6CC2rS7bxO2/eYdvI4AQY6LQM384URjbBbA+hQyfdHnklG3Gm7P
11+x12ZWq6/wpXp6ih+JieDCrujEw3uU0d+2kt0u1p4PVaTpcysSvq+hhdRW6r3/PW3NevXn13wo
S+lpM02nby1yBSSyHbrfUsIfACZYbn4JYMW4PfJF1TQXB9jrEs0eY3GhJwBkbjOu0tqUbcen7h5J
LCgrhSXoywrEzf5Tck7KAH5zuS6V1PwLae1tGIMz5xCdCbqaSHO29Y12FgLFnaOe1Jg6c1cxVLdJ
eryXEOl7wunvmNAFnEli+asNg9xuyxunPlMj5kz5YpkEWoZTJ/BiP/0UkKeFMAx1NQlH3J6XGPz4
MsxITkz1EmjXOctD6yLRWXNIrBTX7d23qq6my5k2OsfpDZWvgY7GNWAQuNp+Y9Np/fbsL2qZuo0l
ypcokXBu/E4RHbQyxA/iYN8a4G8uirf1bpcApSZ7c2Vc5KPkWrsFegj/aY6EQCOFsN3jCWulD+g2
jCVNqYtrIDyVXfPXTufTTeft4DByf3IkTG0kKv3umaXSZn6WW3lC6P/enqjfbgPGk9YDKQJUwcXw
GXOjIaDNd8X1u3EayK5CywrKhYGnNeHUfnKOy9e9RPuA3zXnOSGrlOMe7ZI7M/Nktm/xz1ZtQdV3
EPHdPv3s1K/8+NKd25ZjiB26R4VHNl7Lmj9pZ/eaPWOykGGv0MVcLiV6VP54E9NpImN76V1mdz7v
0s/7PmuR8ncdtIbCweGcQ9Zj3RABPAWVhyU4vPJBpk529IXRLX9pyFQ43Fsexg+PnEQ08YqUweDz
PfE4GFNijQ8iFuV3EEsG/8kHKxbKvGTTOi30CfkKx4L/H8sUokNKhnRMy046qmhAm1LuEvEnPDDN
bLsXeAz9/WHyrbCgL6ii4QoXek/b8ITpt8AydB+WVsaVHjuMYP4/QgYlf2Vnyz8Kw3wkZ2N4jCMX
/377XFwXalAjkFPVlQv2rTgELRx/JbcFwwzL2mixDEizj1q2wzMlLhUwEnYuY96EmxptrUj1F+Ly
4TEN7kzeMmuBerzmicBWEwmKKC6QDAK/+cwO42b2TU2HsEnBzxQPzuQFhXrZQSE8Tjw5Ur2BbUMU
x7t2DxMyonjSw/E7FgwPafyuSxOco3paOdTXEChD5D6CkLmsQmYE+ZLjkg8RelV7qbWpfdq3SZbt
pvKxPnqXseQkt5ZqsEX9OWNJOuJiN1jOLGJRJfcpT2B5nuujK7pUazUgPj/M/VHUycgu/ynkwzv2
2pJE1P6dvpRdMkhCByHyVk8LyQrxAGqXLy8a3Ghjm+Z6r1YIEiVsucRp39bZ894UbzY4TsWro9Kp
uR+S67fEdPZmJMd69MmDtiMaWt/U/c6sAXEAuA61lE2R4SzcpFpvAh1ZvMsX9aBnUztYrLe/4oi8
pwtj+sl1MyRzzieDH3CqAdw922qHDc6VEUUJgiB9hy5MKh+HxkbuoRpxX+c6tT6UtRe0AwZEtACl
I8ia/A1+9TnA1LdSmGgUQKjbMmWNpEcw094kOZe8/V504dlKZbMridSw232+LNzw1+2uH3YiAGfP
F3yR2ejobANeqdqJNZ2ThftYkleWsPpQuZH9yP1yuhU9CY3TYMq8LQJ6oKNv7VO0yG3Zr+em+npD
VcNEr2EsxRbF2GtTtIGlwEAoKPAG03eKAJ6qmN+dOL/CTOHC1SqByi54RAEU7bP3i6feg+KDWo4y
3rSmEPNBnWPYfBjl2ITexl5Z0aWDBil6X8kamRyW2iQ30kUfTChAePNUj0pp/oiefE0sV5/SlyiT
MvSBIV6gBe04gqD+WV+r9v4El8hLHGLtUed/BBby+NwiBZOyZ+bWgDtfPI3w9rL5YB/ALcg+P3td
cJG8TxOVSe9gQNgd780PUg9ubBYIDzoBeZ8xetgL7HW4RvCFptCxWu8GBYFKCgdh+GT3rJu64dn3
YplzG38foti9p/Qp4uflswR4AFtd5TBqdT8UKtH9gg92kurlRghWN7LkSbhhckG6KapIu9CxJSxn
HOuBQkIkq7XSn60AFtQSLGkwTTSZMh9L1pp8AHETqUCf+9oIdJlfdrd9DvQGgoSEPeS9WdTF8aiT
KqBQBQ9Fxlcl94mP7cZJFsL80hiKg31IJqVidpc0Q69E9th3OkewSylitzosFA9ux6dW8Zq0qWXk
ROu897fH5Qn3UNOwlGB785OYIKTJPm7TtguG67C3I3MjN6AKs/5kglRyEsDyOdHPFZHI6q8PYmuZ
c4okdEgAJ5HgP0kF9F2fJUQRFZR2nHqTwnnCUVMhAEKZgu8l3LChEVLsCYG5iXvjQH1fTJOMb8TE
ZNVhLx+UlN0DPl6voxr8t81uql5wGJrd69iDA1787tYXHoZzhLLiz8ExFOBVHQaTqblfnNvkwpum
g3ZYErN1shG7CleCBjpHsHXtMqCX6Jgjxmdrz8oX5eiOjUpMh/HK2apbGM3LFQnZ9SH0IdmKEG97
Zsifgy0lAT2nXfrbs2tUPMs22c+fuu/xHlB7oYYYjSbY6apOidvGoQPLw8hawJyChixmBBKQsBE+
qpvdZr5uXhteGVglaS2ZxhKhFyFi33Y48e+l48LKn7N8bjwSrjs8IHzFlF3JNeaYV02FMc2aPdM4
L+HSEZ7d5oZz5XuWsqffoMVrvSGURsTDElZTcH6rk1yJTlTRtqO4bahQ7yvIZqoFTH/nhFnBQkmV
903hA0qYrdICRHEu3Dk5Eg8X3hvUNqb7aA5lw0h0luX/pvabUcRIxwBo5hu2yhv/8hGb0rAxoE7c
0Y28ju5fmoE3+Ts7u49I5dLPS37UPnCz4aKXPn7KDBT3oZ1M1l/lkHXSA3Yz5sY3dAgBIYizqvsH
j+mOiCAiVTWir/JnzL61cqQGVlGuis/yDw4p9WXRaKUQrJncENEeQLUeiVibwelRubPqLUS9EyLp
es2TjgOk+ATRnASIqUOpqVIzV0skOiRJKCIBiriLJgu7uGzbEiX1uj5XcKlJmE5fjNSL/4h8ZrEQ
66dbG4tOKClqYGLxae3EhanT1+kUDMhzRIElqPJQ1v4h7c/MRS6RJZ8nzzLq/bp48HN7nM8+NZ2G
Tqrs2od3qwTNQzxTKUgZGUK9TM22366kGaSyCJp7ng2kAewH8b68/yC4wT0m+OPNZIWpxTJ7MMQV
ZnCNMUJFPAYRaLadR4W+b+OaSYzF6PVbOTFCgkQsvWrnII4sNMQERGsReZHyeva+3WNDKUjUDCBC
WzO9XU9FAudDm54GXb3zmFzkRt06gGr0yQQkz/qfZWAiB8zxC1f8CwYvDnlzXtQ81xlj0uaXikf7
0E8P3spQevDNtY+sVLWpBoLhzXmGLi+UTC9e2OT7zOd80EXa3eGNURDXX2hduFfoUHiACK5wjtSZ
aSAXWnuMNBOqolnATsGifLlVX3svJT2VrPycqcCb3CEsvCkmEsdH1uNCukJcSEfmy8NMl6S7cB9l
m+mpHWJ36lm/czI6v4p8aRHP2CuNz+EBUiiTgzqOqMN+Tp0fcvSgf3pxRbvGcC4yjuewNGm4qNUM
VVKa7U90BK92Hf7I4jRMj8WFwhCQE6nkhmjnuOT1cg1TlUYP5sj307ibh72QEyacE9WG77GalESd
We4k0JKz/jOwtl5vwDFk6A7syM9PR8WcDsbgD9c94+p+j3llIcnr6fGOMne5ZMIIWnOPULXMbwD9
7WV1TOH6HUUQ4CX6lnecnLk6ZApbnzHrB9P+rxuAcd6LUrvLfEUr6OHXc+oNKSVPmuEcGAeCLmVd
H6NRtTc6WFYKtkFrD3UNXjQwwC2jy9cNd5O42/oSch702MFuRrE8Cl5VK0mILV9ogcafJK3iRyeT
OVaXK2XUQvxmUeLKW4vqdXZ3q7SCSN0g/fo7dK//xJnioRQe7KYEEPb6Bat4k6NoJ6apctojelVh
5uvhYTFDDM7fr+V8iwk+fzu5o0Ll/akrDptkQ6S28cbblONvklNN9j8dSiRZ6wfxsaWwCdpSS0SZ
gEPLUGBMPWd4rWA7IUdKdnoYQZFnUamQ9l8kHvYcIAMvzRWfViu8wIaAoHn3ux3bJI0WtD6aHfTi
NbKY1KuPM7so2mUst1+JhD2/5+QhtH1QpeoMK60rg+y/UunMITUnGp1MltvOAqPNiYdPoqoAji/2
3rcPBLx3HlRmFgiRSMuTf0r5/Da18gHEwLnOwGMXLUejlr6gKfkTqJ/Rkuaw3BBaoYVqjYzdxXvs
Wa3sKSIp7adqprfMACe7+T+grGEEuwkosA9XGCH1DFSW2rT21AV83coSvp8RURpC2k6m/oTlyBKo
lsUV7zPU5epCLLvsknfgVnUgwB1x+opT3B6QDdKKU2d1az7lK/dQga347cczKipAi4EKTy++V1kR
Qpurlon3SgIKEQpwNlMBH9PTS2Irtql0ePq5E48N76t24IRpZaSQhw85i0WSnuB0odZNwlfgpS5L
OZs0vhxLVmtActdQsd6yoXHw4vKyNdNqb28cPlATy49jZyk6npeHT4B1PXElvESEYNkSsUqb2DDJ
2EuV1b11KeQNlqR/5/P1Yk9lUm8ZF1B9aK+Eujc/F0dvxIfGCzdX3EA/KDOCRv7IniooADCoBJWH
XNL7GBbGqFkrjB9Ow+SRjozvrMAhkDPKqmcR0Jv50xmlvs6zUFIiCBfPEwuORfVzfYJVU1S4qDlg
e15BQQ31BIIHSHk5Q5Sz95z0e9ZxouURaZ6CPm0YcEWDCf09prv3/NSGHLm8jcTEz54WgFXdrMmT
ZP2goxVjAHAFQ63hMzLuM1eSt+fCmPwp1Sg9DAcRQzKxKE4WwUb9sF+h7ZIrQOU2yTDQNkh01Fej
VyiWspCprKRHb2WGK6vg+5T/HfNi3VR4s6VKBBjoUJdyV/FH7cMC6oixeWalG46jiCg3JXrNOkj5
QSQKUotu5A2ZdPaaCgOxO4flocr70mfW+YGN0Oef/srKlQ/O2UK4wM++WpxKpb1Ndvb+FaZlrMj9
MlBl6iFdIbkjdxePsf8xlyOh79FPFl0nEjRJO88lpA/J/Pzj6yV1AmRow0jfwuhtbOeTf+CVwdQW
3VYqnJV+kboRSTL3gANu0d4QH8JjduR8TnRpFhsoOMoBt3RJelGX7ZdqYjD/kig1lK6AKsFrxbvx
tT2tN802X5KOcPpaAOK344Y5aax6O39Fsi4pzmuS7bDtl/x/IcEMKE5xNq3kL/HFpMFFxNkh+chc
H8l66JS1j8MsqEpyoof4MtZjSHhRTQ4JDXsP8JbicE/5CvZNDhs5/DGTbRDwL90+mFSybGUZ+01o
Y8rhsaThf4qqYiv7o6Qksvql4XIOlveVHZx25jhmsk3xxyxkkvZVybwNHyb1VJh6iV1EIggtcCKU
M2ZDVgKfsZJczzDlJhlyRDJvs2XrEzJfgeZan+afuAlyPeA9E8oQHAFVn5vX9ccTErmhbCCue4JB
XUav2jOHTAA3wKwCDhe1iovdm/BnAzFYYYXjNs1w2SQmJG+0DspVYo9yalY9rNPXYN2Invc6hGvn
zwf32RF2rJBGJX3KMYcV/6wztH3nOxDes6z88XlJjgwwMkhDhD5E8ikbBM80NVOaYVjFOhxthM53
3BGkSwfbrXWRKw97eMwJ0RZ6oeo/rIj2uXzmfXlRBjpw+2g0NCqcYWhMUpr7TXAi82lrV/NwSnaj
m0tsvSBUnOpKVzav1ix2lFOSElsEMzzyD3bWaqaSZefNhEkDahjPbduoMnYWVn2eBF2MTPqJzW3g
HVR/Y1HMShhHdUqtNGOzpy2rPxKyrP1MY3DKSuwqPONxu8yFv75CySwoHWHyScvIkCqb9aWQStVB
Vp5bKvH7Z3vJDxbojGsIYN3gFB+b6qldjakEtWKxMyomnl+Qtj3+dpFieu8FWz9IpF4I3nWY0Y90
dWuSu3HOiIsa0aNmVlt4H/aj2QJVP0vb9Mw5o9ozIzTYukkS9m9guwEvLjxsp/xb6XFROm08aCki
TSoP+f/Uwz43sqgBXg6rCONlcLujbVlwPgV92KU5GHhjlRYKfjC7HZG6JYqsl29+ayA33p2I7BY/
m3QlNBHUlUgEZqLzwwLrB7AwKVntwBUy6U2PSZ616tihudWRokOw8QtvEe1yaJaUe2YRClhmRbYa
PaWgVA5WGW2BSkC7MhhPkaatnuMx96dGzANXfy18/DIb1S11oABRyFdgFPESoxDg8NLJGKEXcRS8
dWJIwx2t31iGi7VdeQdEj+teYjIKDM4q8oyq7MMbuepaxv87xVvzOOx5nV1na2R4+fcyBVv0IJiq
1LmqA9Yh5F3mUuejn/f9ApOIRI0sRTdXQEvB55tptqUvQO+aqX8i3ZLbikvsA1mC36Ndtvm0OUJj
iJ5AsNoyAYT1y4m61u1Rty1H6EzO0sXVFIaKRpkDnzqA14K9OuW4m56X7FdHiNfKPfREL/DRNmHC
kaki9r7JIeMiAbhfFBajO/cxhszygcKaVzTj3yKnCGDtKrfa5lvaBWnZD0NJFSvl8VQ7bmoQCNQN
Ixo2ur2lijgwHpbhznNib3IYxxcuQNmCf0aXnMW7wzhgBQ8mMLa08HJgYzmonCg76xAOVG92HDKt
slf5xENjbvzSzdMkQuw+2clt1kSLCyKHQpWuKRw0vsSGVYP4wnLuCZJX2wHXeNzl1X9a5Ch+1IQG
hnKVJ/g0kPG6lpfLUasCNoJYWWlivc7C7hSZNP1lqhiSX3ljG14hvjg4JWhZ5mLShlSl0WMRYDja
aH9gyXWdkYYwITcZKwYxjzT3sKhvSZlfeLC1pgvQq9QilTqzSvJpbtE4nX8x7ZjfqL0W1Zk4yUdx
CrjofsCkrTtFMG0IKlTlIWL2jFXkxaFm8ZgX9N82qlMqQ+FcVHiWL853GxRVGfhTUX+l0uLUng7Y
yfOVOcW0AWvJHLMTqvQfWOVx0+3UeXnkrCIxKKyvEnV7y9o5VVwAEm/LnStCmf1Y8EZxA7ybACfE
5qSuiJqZe4aQx6uvotTWPYE4wRolspXAquuITlPIKjhyGRNo0d/YGuSbOob15we7URu9qUF1fnTL
bAMWrDUPG+VRkZSzPGUvMw==
`pragma protect end_protected
