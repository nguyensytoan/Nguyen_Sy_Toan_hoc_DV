// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
1tOdmoym2lzj8IhQOtw2/Oayk+uCWA9XyY84G84VSt2No+lIKsCAbK39CHSZdTasNn+vLfB0O1no
ZgjMBV544FdhAfRyPFkOqIMmYnHG5WKdBYFtAF61Rmor6chH1I0MMppGhwlfBv+cw3USSCensrAC
RToD4gqZrAv8LE1b1IguqRoo96MnZ0cySi2uikpkiYTWp/OE/pW1x4dvghrv3/rv0oICQYwoH/NQ
GBI/8kH2FGGzmTpGIlKP/l7qw6Fspztm2EsxX3DYzIGtegvEb6it50HozZU02RaCSRCsakqpkW22
n7xQDHkpYTs7vNt3+6Op6aZa3f3gjFt12LKjyg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11616)
p8j8sesiFjnNZFtuLJ1/+DhVpOZZOM3kiTVdfIDSaf1CP1CHKM6SFlPRp/EYW6KNm+5kqDLeT0yO
kd6GYFYmPHTjLO3yE/vX+0Z/fOlmrJ6JkB7PInkh30Clq8CL4kYucTLX6OtUaUcrLYAuQzOG9mo+
HoJpblRm7ZfuxREw0+RnHG/MF5rvqNIL2Ofz8FNqysXIF1WYVj55Y34wNoKU4XbGrPms7NJTj1Oe
yr2GZSxFjdhvEikwl/Pr1xsf3EnZ7tpeMNqPVUYaJf0O6Z7PFEmmPyEaZh3QlAWI1LV09W7Grox4
ms1CIIiLPhyKd3hAaKLJvZG/BGkvVOU/cSMdYSvR0pma0p4nwunIyT6Xh0LyZBK4rZ1pmLuquYSZ
5tLyqW7tQQtO0405PsgBjMe68uXCZGKAdl3UCOnc+voJIeIzGtqa2SK+P5i3do2yS4wazlznaUdl
xvGVUCZiIpR6mGB4KbZL9iSadYbBIt+b+0Lex4mwSmeChZJjAFpXzcD3/r/QG1S5MTiPVI6XHu5J
ooQbZ77sTddbGwSq08VHqAT1lHKQbVYCDv/vUkz8nuo05CQowmpYrIw/KFd0Y8i8fAx41ysZtQ0y
8++RZ8YGguRTCxAEi2QU9ZpYASi0kbrEfjaUgUFOEKlvTplF0iYa+BNVq6B8sIBUr7W5XPiTFqNc
3c0zRo/WLvxiis50iW/k0ljGov/YJXDp0vpjyuLcg2iSsXEFc6N1l8dw+0tifSPrpgaaTdy8plS0
cD07UvXaYH7D1IpNRt0SdrH6+8gRpRQRTGSGl2aHjhImc3FIWlMvjdXil2NVIEglFIvr7BHWic08
AtiJ0UHCoercwRQlOBeRfTofNRTI9U7xKzPolbT1GzkKf2D7tQQorAcrULvjqWblYPZ+9DjSDpxx
HVMQSyy4OCJs45IWoPXBw9K2HFu8aDFZ5DvQzdWebpiYfDfqBKXJYXZO7KtGlvvyFr/dT1JijhJu
D3agWbgwJ/vWI0/tldOFH8la4CNOprhzyg7XINma1E7jnZGDrSdvG/WH3Dy3knb7EEr9n+d/GqoZ
oyiPqUseSruzdWLwMbFAdDGbDcFxg0lM13eNIFXquPPsouCOtuvnE+IJiE76CVVNegzjKz9E9x7Q
+t7BzaxdGnlqBpTAR3vy6Abn76ESdj++eY70Xc63J+9N7pEHVwqWlmOjpozLy/NsheDPB03ldBDD
6fxxkLdeGLh9bn5pz3zhxBqlgn9DQh2/6OrLFmKmsIby2K41ujLG9ovzP0k2+/C2xuHrvDxzP3vJ
Siyo9Ynis7WZ2iEXrzrLZOOf2HS89G7rZXvIgQZy6M/FfUt9KmhuMf4nb6K013RRnulmd6kp5m03
cWOeF1byjP7PigcG85KllAE4r4uE240gDqv8epTHdnX6uZRJaO6vJ5lohnI1KGVHzvqmzmCsdkWO
MZ/HR/zM2Ql2/E723PjTdXRPCt/Qbc1wkhruopZllRvJ8BTnMyJuDcVubtbBKgaoF9Dz+/aCwFY6
gH7el3JGwjuQ4v/crzysuQIk6f9adTW+u89U8E+N87KAkoYTYkgC9yeNiYdusOb733EkAMzeb+d+
+m8jcQtsGLzcDWGYhStBwITC4LXCEoNcz3ZjyIucmP1SUdmS6ehehpD+zY//U5bjWcFrvH9e7egf
6IA66b7Sys57+gVzvDVMN38ar+f1Zv9Eynq0MMK9m1Mz461iDsyUGREH2Py3YsN/fF8MywGuuGnC
P4mVQvboXQ7qhLxBcu+X/GVSzbzhKEANqkpbmYeUcYWUfPofKAJiYz7bNaLoWjuzPPFepDnXVNuc
JrWu1qYaUdV51DmEh5/wkDPeWq6Gv6uXlBZQ6f+RcP6YXJ5Y5xP82JHYbvuQpTxkvfS6bbwyBjC8
b9Tba9l0RZzeXb55yk6jmTC59mz8cJaKHiBF0w40yYVSFvCRxrb+c7/6hNd80wy7dYp+T09fGTpE
x7gumeHtv8HMfifFe9YfRK2A0EKKs1bI8D5IyyUFebQhy12+ttyr3UXetAh3YDhQsr3OVx4ToL+8
ooFIscNfdjAaHVbJlapgsBhmezn224MPjBQ2hb3/Nub3jQU6hnXooKdbkdR74xyH5KMpprsoZz+s
KuxZBHfK4YjmUWPlUYX9tyb6P2hZMGgSOATHl20b+iidTDZ7/1lQlR4pQKeAeXK1gecvInEbyE9P
trgIyBRmiUd6kW+4S2wCk88LwpgxZh1tJxuT3pQijM47irKNrgXEH42YfJP0V9ORjGvH+HM4h2DT
fkuiDFxoIXo+VZtMLHOaI9/kjZaaiwacmlsgE5FWx5B7v3HkmLiAUNN1nQtOAb4aGa5ifT48mq1m
FMSbZ6cdGBKRLoRpoQL1r7EawLzh9c32Dw2tM7Ht9o+LM3XnuQUNBTx+Pa0jl6xex0TwXtMQKwCH
3UAOFvh8NnayMZY4s3FH5FRXZwZtaNsOOL5kkCKkcPVDGet6J/l7pXd4OkhCg0hQEi7dh2qINtZ/
VErUpfDryepGSnQZNHchPdAXgaaugfXh9vmXORmzCwvnZWrmdF9GOJtpGK5ja50D/UUxXJCq3rRd
rRvMGP6JDPTW5MSLYIMC/J4k/2JoGG0WsW0ve4usLl9iCVwMUE2bgqBpIsrvOS71ZVcQsLT+rU2A
cy8GfBcBrcmomDTij2S5xoxOoXhg9WLZE3HyVRxhtYRWVEnICrjhLIjw2pZerDZ/pdofBdggyCzx
ijWOINC7dnBy4k3GBT1QmYcpLKGmzaAZQ4nvleId0hA4vgXrVEczzcF7k/435sQ4QDX17Lx5WCMv
TtFNAxA9bKHkLVbfCyxq/7YhpJc1rNqJpuO1vxWoqnfkmIzRqYgIjNgkIzN1LA2Ybb7A2nH/KsqN
lTV+jpMOaf8N8bC+SuALG1Bftc8hompbnLKgHqr1P1wpY++l/KiNS9fyVfo4Jvz/pUcPANezj3Jn
zrnXWTTZvkrNriJbgz3tZZJD1stR3zkl7M/dLNML5yBu8yCdqIGQK0cEfuMQyDS7F3gyZUi5IQPe
iuSdzNue1V1xmTew+pO6h0Ph22E9jxr+MXzBOSBsgcCFKewEByM7SC6PVMTdfnSOkbDReqxUMpn3
FU1lfBmU0C/9LkgXCXDEWDhUxXoNutnAQdYN1YZTDr7M3eNF33rt8+T52dtQIptJc1eOQlCrYQ8e
uw4FUs8UYbIMGjvRKy1mZO5pNEKfEFB+oB22rceKnPdmCZzqMxJUEZrRifwg9ReO4ks+yufsyUXL
jtXyrBZ92NuPKo1FVbV9EM0Gu0Z2+1AY5CUhqRBOaLUfeQlFnxp+E3+6NyzuUalWxFuDzLD6JOHf
duta5KTiFeHyGDFktvw8IeMpqqkz1jncCt4hl33JU3WWmipMn+9vKW0s8RdNO/cBlVBQ9RK3Lkua
uY7iwiqKd12y2yUEDp7yPkK31oS0k+4k77yL7GFiVnGSUIGWY5jgKNtALOVH0SC+vVSB4p9Rg4QN
80Cc/ATEkqaCzKl6EyW8stAbN/zMR1ZPwLDq3sdaqRZfhvTxv+P5UcyOfIBp8XMsIZhn2j1xLewq
aBZXVdfoZewKWfvTUvflPlVcUhKzjmlXyNIlC0T/XLOsa6b+SYTvSZh9ABWVAx0tigut6b0MUJCW
rXXccJGj5MEX5YxGm7IkjXvzIsV/ZACe91VOXLZ4/JsFsAUc1Hsl+0hluDk1F6kxmG5/jKilTiXR
al2/BZ08h0dqPM2/IQGPIGOFMKKqtfDdd6fS5+5BcOEF3mEaQYDXgaXvoXvfsnzv+hc3BBXvRTJo
F8qeph3VjR2SWVd6IsZZN1O7IbEN/vrOZBzUCdvqEDmdcLm1VvaiCisWPzVcKvomREqXBiC6T52p
Drfa+pwilvdl/KEE1XHvG4KZzps3Ok/syKHpIFGFE3eoRyOZL9zp3aEsi0ZENjJ3hVumxZN0oJyE
oYy1INOIbLQgcrpUPP8G7cKOecu2PT8kaMKdMIoIeGpr4V/pnq/ALqmLjLvsujDhNORA4LbVKJpG
Pk8aKHLoVRiSEkAUtzLQeipbaMgJafVovoMfTsaUeXMvbsCWaok/lC+Dihrh853+dCUc9mg/bLRu
SJ43gSz9xXaAbLg9b5ZfeoCcl6GfxnkwtSs9PPfDx8/oQfEo3i2B5QA77ljxKGf4GAIHh5fZ8gXO
IenLssl/WU/h3TdM8TpZlnMTPWiwDsxxK//6btVtFYG75up0C12ncNWlgTdVObZMQMA83G+qWlGB
0y9+AGVyBukIGeKdaCEXyxrBbR34bYmhgTAHBbZ0Dk/4S+n7PkxXJYrQmJ4ghuWM+EE7XMAidgVS
P1Tf99PlPFm2xngnD/0sTeEHemhGEKidjOO3l4yM9EyZ2r8hCLm2U535VC+ThstqpDQc1n7bnkuE
/ZsdzDY9Fk2HoikNgliqm/Pt0zV8QuTqICYdRDKHVeJbkEAl0IM2kIsuQK8kcmyGXVU9MuaWjupd
WNb1qYxq3nlaFnksW+3H8l3lHlqYhfWsYTmuk+cQHVwA2u5q4jmGpjXbBjrbZy85DlaFl3f5G2Er
xtQvkPdRN4mefHG4wLm8HWbJALu5AG4OvnE6Dt7QTGsHoZlGkD941zP+E9AX3Iw2LkY4zy12Zi09
wwpHtuJmMi0ZYfHrtjNUVXqsbOEXtgao5J9lw/WYzuWCpqOmt/0nAqvyC44t9OvHLcCkIM3nJhOO
OneSoiwrJxmXXJgucsuznL4Ofw6RDIndlCWJIssqAdY1TbJQef7MHsZPkIhGQ6SvqCDOCzsHScrt
6nC+tnJazNg9LHORC6zgPl0lzvWIAb+yzm1S9mq462W0Z1MnicPeEORkIYIu/d7BHNBlyWNyFLCY
hMOsvsv/eW5oyO7vdRwJzYVPGOvlhY4h/Hh/T/TXE4WOZUkAT3HmM+fmPy26hSUpLJw7+4OnbQPJ
pF6z8O9UIRKVjGq06PIkP7X81NkV9Z1GvnjzcvGVtvG4p0bjn4bMSIzYS3YfCkehSkxDf1eoIg27
rqOFLJ4FaItPGz0XiJn0n8wmJ9Uhwt4vz9c6FXQ5K8HUdp3zASt8jKjx2aUREw//yIbEkx7XJVLu
/AAD0FArKqLlFQkDlscRNvdCPIKCZNqNrI1X5gN+fIXNA5C8aQMO8jm/cZKtS9rlCLfz57HfCtVb
aomAgOt6lYZ5bYX8/5P7Q6rBEWyGAZxhvwaP52J8f0H9Ev7ZY4RZrBRq/dxsYwfbHflDc2TCfFth
1f9AIZryo9T0rIJqt5brWdpYLfbhEaxka9a0CAbt8l6sUIV5ofu0+rs9CBr76TgOQlwZd97cFo+o
oMb/GZyfrnBYYpf9GfQ65BkTG9UMm7XxPWUF+mvramog+4UOpbmTSuB3wFm9GzoNZPoHj1PX7bH/
EVSt6vZM/kA0fX6sX5/IrWCHndjJtUCd0ERqchhaK6JlHyhPSuhEz4e8NsVdAOp5eGje9cPfnTkx
SycBJ05f3jE9SBugxlBzRas/yGwzTzrWjbbrdvWuNoRvhocCHWvgfdrMjJsjFkJDyJWo4qWDzf3t
egPLpPV4c62hUKWzFQ2ByqKhj6g9tqNHzCi3V2sVxcSwcNhy/Is4HSE94tuwau4af/lmcu+WqopR
4oUoONNFvo4i8Eu/GSBoy+U71+cEvtIcxPYLW+iYNZwUylMmsWP1SL5DamMZ06bfRNTWVlpaubWc
YwzxlVNBwn3kVmICE2hNKsnLuIBLoq3XKewT/6WS3Y6qBVy7q8woW43LRlY2mJDcU+lf5+pkFqYK
vN7l+XpQ97VPwwYX1a/T5BqtRIzzI0Jh0TksD6/eAvWDH4A93Gwf4eiWQ+QpBq7R0/N6i3GcfyX3
iY6tJkVW8H9v6i4+NqVOlRQyyvu1hLQh84/BUDAgxa6vlh8CZgiSZaegM2jgKzVk5z4sAQ+XYpG0
qDc1Frfz17+4aHTwReB8lDSjtJDuqwtrUpigbBX70eaMQulqyLxjxzgnnHcJQmqPWOPO+TzIdKIu
gwOFlSqdMc20TTrJRLk2kWRwqynRh9QleNMVfaQHfIupxmc4SAJE/NE2PkGexEjL3T9QhhIQufyf
BXyu+81qyQxOqD3UkjEPBCYZiOmMdNj9GOzOKK6lK4Smklxmqv8l6Tegl4hQyfFhtnkgotKY+tII
dGojaeXSf9aBMJDZdjYGCmQhHxqfI2bqARxw9SpsQmnia2mP6pARVHWx8lMuYzTqAsb0/3+kw7TR
lNUl+g2MhUSUpF7nSl+rZJ079XlGrxr/XuehWrb5IEL6RwMrq9etzfTI7HbTejwh29OzZ0Rhrd2a
584CQIMTYrWjaJRSXYfSLN4KAKwUTkEs0xvjjN5EFF78ZmNVf8Je/WKdClPa+2UWfd2kbgQyMgX2
gSlCOD1FMjL6lEVKN/H6H19/CabwvAI6lfDMQn5BB2FC7urN0yUJsZkAIs4/fH8WdVPI0NWdd1xT
6gW8IBItJsvDR+qstg+fD/tZWFPHgD+CcKod152yGzkqMZlcaRdT3nhN9JECxOzYX9R33baueaHT
aBKHyqCAwAO5U5QSEnS+3UZteTxVzBzV1xxnSiror8ybeGayPGvdvQbEw+wt0oM2UfV3L1sFg1uC
ntPhYZJA3t+bsqLHgkNKVWmx/ImjnI1TGY82wNAcanKWLOnw+CoWU7UvGgVrRLvm4DLcf8bHH4nN
WHLTVERCVjZaN5/TghNdvbZnvJA6cJqLs/2SK2P2oFBSwbyy91trDoqbWGpqBNjlR7Js5Y+fpIQo
EzooPLeuU8P/I+hNkwRzRQs0EtDt90ZC2rsvj2t91t6U9RD7TPGBPrl/CXmaX2mf6jp/WmCHODZk
ezkRCZmbQkcT4uIQNXq9EaVnEKNzIVqXxiwGOjNN9OMXXWpWzbPVES4vFMkXofheyjj3BBhB9MGv
TYu4BU/WVXbK0CdCkVGDnzuuFA5RrdShTawKoRaqyUSEHz6IODjRHT3G25vSDIdce26bKFmM9zVD
q5JruvKBcCPxPQ+Ytl55nEXw7lvRKjMOMUStL0JSex7emeeN59NeomZIa+mQ46/PhVSvA3HjaZwQ
et8wx8u9j8lU0Y2mF+b3GbfG724XQcjIp67SH+3sH0dV0dMHkkEy31t3swq63GCk2sT0oRDGdrFZ
r+7JHjef6rGOiZdS9GNKm/OYAcisVEmkZOly7mHfb2ZqhIYCIsgSJtdFdPm9thfjoXFov5GHDX8P
4VUVamooWEVmkp3UzKxci2qxkwSkmlWC1Y+o5EjTE3P51cNlu89bazUpkitfq3HbpD1aV4UsJK8F
fPw8pAVJmujku6e+C6Cm9cNtHxcj/+LU2ajFph7GNEW9+xrBea9bTAYL5hSMXS7jp94jp5G4rHq2
EabFr45VGMxEJlZaLL3IW6hqinXt+BIVitMjFgY8D3Ohdo0IdDQktF5ogZCsviuLiFxfJHjtm08B
/xxX5LMvx+aLcQgEudOC0pO5b95X+OLjInFTSIxWeqV5Wg6V+5H/pjHKTLcXl33IkjYaRSdhAB/h
4XL4ihEm/SfWdD8tgsciSM8PQ6W6rUXmenoqFxzZq27WI0Cb4XwRWk4fxF3V/pOIdjDKQEg+5ebQ
76F+wGa1MB6tNlgMKTnyzMcSwDDOQ6T8cosesSTVWSzqQ/rWBD5xT21haA9BtPVUKuMIVyrDyzAA
MHQePhS/QgzvWaUYbZ5CcHXhVepQENUyvWDySeWH6w2r/UEXBrZIhqV72rhDxoUGwcdpYmtFa1Sz
WQIVzFjUaXfmBfzdyQMB0vW0z4W0xvhtLJy/VGGaQRuMTd4ZzHDPAhR6ODLXQvHgwPkCGIQ7zLQ6
oM/79ysa8UJ3J4XJT1GF/u4yl1RzPMXaHtoR6OJ8Ag/YP1J4RmDkeaGIYpQWHe/j4r6w6qGyJcx/
meWYzep3A/3S1OPtWAu8a8V4eVv+dWy+yLFYrOd751dUmtcfZwjkeSd6RN/GrCf/r/xXyC5cyEnO
5Ou7KeOTqtCjb9fn05ijkybL5wczpChWzR46Le8nN5Mmc4W2eTcreXFy+FVqUvH35nja1IDnRWwm
dtHJWb9e+mCRrtHDBZTwv6WmwmrBqY+4q6VtjKVhFoIv/B+JJzIAyopQxGR9WmZ05k+DKj6UajyF
PCr05eaBDRrtyfn8A7NV++Z7LPnwE98Njzdr2gruiCJa1+rq5d3N6b9TsA8iDBy/GHdEaoWwP4/H
0ygeHnL3dHK3335xuER8mebVjIPRHAPivW4i8dQdKl+3nvV2bzCM+zobytkqFFSpmyiGDuVbwMV+
gv41Ro+FMNYyK6s7LiCqsZF8FbYMbQBGIkd3YG5VOMQ6odlaSPxK7Nnht7bAQk91NloKUJAzmhbv
jxqTVZuG3YLZon1HcZyoPAmU/XtAzLodhy+BKRoK0NtggFEh8U+pk8S3sK4jwQEgaDKgIjVtBMZu
Nk77Y+F7QzZ/UrXeS5Dx7cB/QRrWyVAAQNilV9IR1IRiTn8tJ++G10kl11g0aCRxMI8B7JPwIw68
RWnrTXgBA3a5L9OZrOVl516uI6ukVuPdABi1BXHxcy/kq2SYY8FcqC4Jsa92WQU1j66c5HIL2zD2
OdsadiCfjigQU0yiOclDu+ssDmXEOA52/mYIJvTAmV/mDeq9aX1DUEqtRG5vv6d+y0ds23qB8EKk
Vqaq2Y4N9TyYnrrz51zs8x/LKt8q1OytITzv7AX+9uxy8K/3Zp2KGqTLMuZxUK0YyV13DVkt7O8r
ZnCgMzFDnOcKfs7H4k3Cf7hiO6IxFrVe01U/Wp02rkggORoVHAKQAwFthfdZE55WBYc3DhYSRL8W
+c3dkHcaSLGxeuXdrxJ4dT3xChyvsq2M5RNnDCFiFCpn2RVP5X66q/N/dVx2MJZES1xh2zmHzB+t
ja3MMBC1zJL2dFGuROX4jFfaAFJascVic01ABRKfV7Wx37dektn+/3ZlBe57AltRIkWWO9MNdYNJ
XtWqKnUO5scf0j1B874Fh98jEEbsX5YEgLx9I8XuQjvERWTEtgGVuPafi2vYFqHiTB9iCVnHADee
J5iXEYalaUjNxlc7ByCe00FXFtR1FtMmf5SPrGvLN/J7/UZpgwB4Co+Cce+hRIpy67H7IOKBSmg8
VZJGW0LEwkx/o3gWwmQmI2RNXWiaCI+XDtDqSNRUrXZT25m7MZfaxW7wr8WCQg4UmNM80+MzlPs5
/GEm8HQMbn124spC4E6PDQw5zj+VctVV6dnhka6xZBcgaZDqrQlgutg4DE/tmFKDWP9pYkjSEojO
Gmm7KZZAILYmnMw3VY5z9YIS/mtUZcKn/VDSw7Ib43FojKf3JqAlUUGEUMm0gldKMkJ7bJyivbjN
MyiEOsQpZWd7t7gK+4BBWphFKqCEd7VsSkhlNIDuGG+p+EfWBwhVboqcM4UTnyXn+aZXipS0zikD
yCNwXw2vQKauGGUAabTgcSmpfVgPfJS6Kky8QR4Rm/15H/eH120eo/YepgKo9csls+TFa9bLjDlx
KFV/tA0pwjbPrCm9NNFon/+BGV31Mk+XVLMnNJQs0FcnCU89v8GSzbQYGXKbvRL6txdqwQmi05fi
1vPjH56xpxZJL8ltgQx8wzDkps8b6AKwBZXcWDuKFa16+zsZJmzCToLBKTFb2/zxcMZlIYL2oVMP
6D0dnbaOjYF8hkMvOAH4Cnl5NJAkKdg3kKH6AJ6kDJY+HUhtju6kotMMjiGQgvlHuh+AVkskK3dz
8iuxp/sDj8IF+QnVEhSARg3oS+qronng+JcYhWTbJ5p1cNImUDeIw98eXQmvTeAICPe5O59OkGJC
v1mToFBVAGnFvnfWaEgNgePkNo8y1vml079Mn43QV3pqI6gtB4El74xntp1kxtEDZ3JALKbezvq3
iv5M+hYlEpEMtQJYqcAWOGgWR7z6A5IpMCMXqUQAP6vd5Idbj+szXEHSw7JVEwpEs3qcWCB9TrAr
1kETPfBdAcXkkDp3pSDg0p619Nn0cHkLFCpiqUdWnzTaKpcLhANL6ua8oTC8Zt9aq8O0rqJm0Uo4
2xEDBZH3VYVnHfR0e5qXpu9wyl1VXOwchtaK4bILjHVH/gxsFprUF3EmupN+RB1mecSv5N+cwo+3
DIFEd18IbBZKDn+UtE9BTbCH2vtwxkyxNWMmx6EssTGp/oyIaYVMryrs4ByQRivmwbyOx2DKFWFQ
4GDyNvvW74YsmLdTnVtGUhc8LSfLBnacyKgPrUc4aN1fmE7kIRzJq/bxiGP785Qgu1m9WXf7RWeQ
zWqYNzqiDxOOzdW1MrwY4QZ+78rIab4jJZwwnGCBqJKUJncGEoN7FSzZZX96RYElYBHtVQUbR/6s
qSHWUWeiZP8I8J4FySWIRn2FNMxCGru088f3NTCcoWXJHWp0Sg2mcz93DCAI4qOBJZHP2VRGWdJK
8Sxc+OsEwBqfLtNOeJWezf7atjk5QHEKcPlmK6+HgdEny3gNwWXGv6nMcvf2KbK2nfvvd4Yx0Wsl
YXqu0J3JSs2Q+9iw6JWZzmuHuYfze2ajBE7lzr+u0nHMt0nUAwqc1hQiKsOS5KZuMRba0m7bSAYE
WOSNYoyg8JW8yhzRGcVW8l3lqon7SZ6zzzL1a0tvMWqmUXG+016c5iAnHIiecD2STw1hyTYOnqXi
3Tlv76KMeCz8AdTZh4P8WQuYxHdDFWuMrRqjyz+pE7Kbk+8okrYeWTw7nH5+KiAom1IbVnqpSoBx
mXoI/cWeYlP0iYzCxkvPujZ3yipWQnperG1UKmUc8b1jqDLShMCZc4cllB5pLR/nrQF+C6MGyA+I
fitTkoFGG5iK6lkrbl2mJWaHA9zTA+yfCYHwRowgB8VVPijcAJZyreU7MfzxikUKiruFXOHnGmOV
UdQ98p8NAHhYEFzurScVRlSPYekmB+0CJ/MFmEkrXqiQMX2m8X6qvIL1PkR1TdejBYJTf0sEVHHe
sP6jjFkBvgiJbPpKC2INdZXncGIj5Y8LEOKjgU9dMKsYsPSGg5Utv3LsZg6HMqujJScZjH1WUSVq
wGZvvRrHRtK5BJtUv4oOkjB1RMqKgtSdAbI6OxrWoaH5mY3R7aQ7wE7JqIn+ZxAyLQz9yTebANoU
rknaGfJgMMHFaTZixW8JxJr0YI7akcekFhgT+iQ2leuWecwg7W+G1nAvySgQjkW9FvKaoPkf9opr
qyxWTKCaQDTnufBRiZeYQ/aL5zH5g+ubZJlZ9m8dLlJhaFMPHIZaKoyuZ+raCSnuGD05ajvWzZjI
XQuB/Z3Yv3wa626p4Ak9aePXoYAnFHn8DGaxwlpo6eLyzleTbZ/OxjDHDPp2ebuYxlJeBBDflypC
z5hgr41sZu3SewcduZnLo8q+51Byzb1AQ9JQBRnhN2xnDD7e5BsxXik4fW/C4j3eGzLdFtLPToMR
eLwZGL923rINX4Dzkiju8nLo3wjJJc6CL5bIfBKAEPOa9v36R4uWhtILqYnlo/k8e2o6O6MA6VoI
liNMPyVcS4KfURmRVG929pD/w5MNQuroK6HiyywsLWRLshZNSUpeeuWNIlDINUC9qvCiwOgTJ/bk
GJbBJ6F9E2fOueSwRjdmeOJ4YMq6lJhixA2tnXWVIZTd1aaHi550P0GGZJXWuG3QdTOTw8Rw2HYb
+G5F1Ewci8H3oHpOIZFkGwE25QhsIZ5kNu1ytUsRlkMzeyKJGTzpOzzdGhA6CG9mZzF6xqTY5Haz
Fz6QVP+NAyUXuSHtV5cu2V/zxvW3r9TO7xMBpVz9jjZZ6sYSt2gySmSNntK++8pE0ExqCFZkuz+h
+ooeLAC3vcLAgJr0P3DLxMJobJ8cv3MWi2iHLyOeeANFKWyFgpAVgW8LkEELn3EICurIIlZkHsGE
68Fb3mC5Bk3aOfg6AtmKwZx2nIuQfvE0sC5alEJs+Css1WJhq+ra8yzi6BQHH7EeCvDLHEDV+Be/
gwzFc4ymEMWEqJ/U2CqHNzQY5MPVFGo/2LFJw5hpQgKYX3Vn4ccBP3hALAastrzznVPOz8n5XKvp
4+0Kh6alKJ6CHqlI++q10pPwBOcAh5PQmqg03ylr7ExSFjfjB9v/pzskrbbkRfcsFfyI4O2Zcv9k
dIUjpCKcpDAzUe+Le8pFghakyB7tPHiVr8v4a8JHM9cLjL0Noiw9aYh2khWb9ZN3cpUh9vqErnxb
u/YlTEhqx6uBatKPFMD8jJ6vMQ+h4JolBW5x3SoRH/YhtI6JrzXYAGbEPX0SudXzJsg9O20oTvrl
9m2hFT/K7Qzf43BSbOi/tJ1JHyNGvZO1HJk+nuQTSSZGUiDYdskOMxmMPIEaGs0L9pLUWDVEvSbJ
OgcVp2vRPd6DUXxtCJw6RUb0xg4RPOSRALj8JkAF0RBLTWT6zLiPwCd5OFhVkKTYt030+RqxJWwz
E4ogsWnQAE5NPcAZilre002G+s4xzJZz6XzM/8H6Wnbi6x/54bGL4rY118EjPRQ6ac0R0sZiui1p
Pm4S+t4FqR3cMFgJysMqzI78olwv6ehAiawLZEfMJ/eUMsatdI6gHDxSEUNDxBZ7357E5WY7EOdd
ncZeQ3fHgCQkZepRfgneEUVNVsYSaYTAeioZ8tcOg5mVFdfgf4K5XwlErg6PsyktmWf/bXSCGOyh
Tw6K2PnSvjOQKlXDHVuI/DRqV22aGIuGpQF7BbtflNENi89R26yVwIBWPSSCE8T7JcyeYwUkhABt
yDxq1Rgw/Jd179xQBMP700lPJgl6KEuIbYSSlKSKVOVpReeQ4On34HxAroIotOr47ZrxxdS16Uy2
sA1x/Rj/MqimUZ2SJRUTJL6H/6hNrhHtI7KKPWyzSv3i8INKhBTbOFhKGLxkcDmMb1ZbH3ZVJa1o
1ZMuAMovo+1X4VY+Wii25aB0dsRq3sXpGrNGI+nI4J94F3rr3+cDVVnd41SslOSx5wIa0teX07yM
Gt+3OxyPBGsN8Ps9f+YL+tUDqyT52G9erC7jadgkKPb2tf8y4e7l4Z1uDIBwkWH3Ugsp00hXoB61
MlpvbNj/z0kVXErR2lOO5gCFJrExTsequnCvfrJMmnHm29JMgXN0pyL6p0wHOzSuxX6MgQ9G1upA
TOkb+2Kuegq74G9OXUdyEqjkaxcuKMXe5Z8W9v0mRJ4zxnfiyUcMXuv8oxUH9mZoU9l7BZyxoiJb
lRlR3C1VIj3HzTn3uMcSiVvR4s4NsRBBJXxgS9ODp4j4X309BIVBgiAjqPmS3mAaqz1io2MmCCl8
iUGRUjJu7seiQFOSUN2RO/dxFEkKqmQIP1P4dsQ/lXppglWZgS6tEecDg5MOnRHEVCdxKsUB60w/
Of+Qs3YAlCvtIXJvKsctTU/V0nhaSeamxQ7zcdWY9K+DYiYNXykUK+KJX/KnJLhn2YJdeBi+vNvY
wQrOEZ5z7+10qxwtW0D8bMAuKjBSLmppR/Kb8T12BUxEX2xhG4F97oFUH3Xopq+d6UzZlwHMfUxw
SO0Vbt3BXeGNpEDx50eoIDrsUYfxKYq8loG+hPk8oYcqKvHWvFedqJ04M+zqYoyD4MGC049jqww3
aYoqPbpsgg2DbIYYgF1AZAPxigB2ZPiV7FKqX2/ehxGdVrGJnjzH29OYVgr/KgBHb0amfyp6EB5E
DpyFuJQa2GPa+Zp8NwBNdWuUlI0MO4STDsiLQ6ZuZ8LvSstDLd1VKCK5SwG4l2/W24dsip/Gfr6S
uEhpqy8wWkiYs/VM69hxcv85QuFwo+ZBMBlH+vArcI98eVjIcmSvq5YFF0ZGsjPQXm7XLOJsyXC5
FdQHgevMQqz4p+CDRDuFIYXm9ue5elLXUy5xni6+QLGt7XVPIfjqhAM+7BHeZD/DJLBNL/Dwox5P
ys+WTELeor9vv6bYkfVppTI9kUk0zCw9ae2N5RuFM6IhWyDPYroUP87XFXm78eMs7bKMrBVe1U+X
fqUl/5Bjghn9vaoEDQ1gxQpUWePa6cWf4IrBAfgaLzv6l7Qz7aiqthWsZ1qbv8OxvYTSVAFPW3uy
cliy/27l/z7BsZU2zEZ2UhMzA67TkPYjLLxm9Qf3biXLkyzw1aJwaI+oRS9gcmhslwGQEf4115Wd
figsIHwyot0COygSh4Wfk+bhZhrIAjzi/zmzcPcnGkumK3WmInAfcFOrHC1LgzaUmqPnLy/Sr+ka
uCeDCwa/Ht0pVsQgybd05ToAcUVoiEQc5S7wDaBTBXNa8beI45sVvGUYkDP5HWwIl5N+fgVcjwO+
x5hCufx/D6jfi/6/NKB+d71G0TXI2JWIKOlFpjTuBB7I9aMAt1VH6fdj9gEqhb4+RPlvYbIzxQVC
LeRoLQctAvyOs/2DohfaPBsT2A1DVYo4xp/ksDLQ9uENPgeuv5yTZNq2mLmLNUwZ5va+StXa98d3
7KwvTizC8LT/vT6UvwT7dzwNI1F5imbTvZB2qkx43aCHFKx+jplOKSThImQnOOrhXk0YFJeRqU9Y
EWu5kUfE/ErckDkIR/RgxEK8jmxW6sPXDN3PvmqheklWNjmRzCKHj2I/n2yx8dUiqFyedrUPRQ6R
qBucLkEHRzRkaMFVHd8o8jCDQA/MieI8RaT/+jAoV+c3BlBCHGMFYrEe078uOPN9thsSj5AVajMy
O6ZFuIcrAAt9Lnpe0u2xj9dk3xzzjb112/dFPsjrdJ/VvWm92IJGIB/X+CbR/nShl4rKOXeV7EnL
GKEIPtXtvFqGQhVXeUCYO5wE+yOg/VBAkv2ZXtsFodIb+DKfRkZ2k5RWV6xhh8fQvItX7eYlI3BW
l9+/BoVMGweJgWQVaoyxEG2fvdif6E53fZJ3Cfd98ZpxjLl/auX+R/01kIEP92Sb4RnWBNjLWwSf
ROSjuSTr7p5vCclfOQSvx6kcdBQz0ig94FNX4OYzC/r4yOPNhb3R5XyaQbTH0Yh6l8cVDmSXLlc7
Hg47Pn+ygkyKPuViEj8y1xXL299D7Tcv76h3uAkq5Hz2yTYWsjfxP5o6jmFB+bybjowzpTaJ+gE5
W0k+v+KeX8LCYm/RIMNoLZzfAnlqHNMOcWjyMR4Z0CQc9tNFfVALEmW/fRfefv6JMY/WCZ+9XbSW
l5KYX16G3o+ZUIAmSoTu2KrIgVkkqv2lMrZsHrJewHf6AOE6KcwJPxpuwAlAZrAS0AALqJKBtdRJ
fIU0oZ2c7MZJzh6xWSWsn5aaBJC4fdQpEUNYaP0qCef2C6MPjk/Pna5GjgbCf/dKSxDSji1YXqJp
Ih111+sy0wo4xQXNtpyopxkGgfiP0LIUM3iIKaS5hUPudWW9WqMQaWBnz5B/MF6sGQ0p4lT0gbWx
/F4Pl9W+YluDFa5YrfeurRiq2XmG17WE0HfXaZYHLIt0+n1DcRqZWKGeHvBETMKZjJjMIAjn2S79
jsIPoRtRbfQjwKCf1sofF4k3DlAEY+J9dAOrQY0vpyIMjt5TN7VDNQHgz2ack/1iOIgPpgdULFli
qi6kl6gJHd7aP6o2qCZ+Lu0t3PsAnJChKEu/oZpX39sTA+7qt7thvwT9rlq6
`pragma protect end_protected
