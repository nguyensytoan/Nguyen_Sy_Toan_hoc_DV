// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:32:02 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qAj4v26jY72kYvD6uZKhN7sWEXx9kkFnDEQKsGhj9Kuwl3K/6pqcAOyWPZdKC+7P
i7eVPIs6vcbW322ESpN4PblV0BSMFRuC2Frl5sahPVG1IBn1Q86KWTB2WFThl4b6
RUaetMvbzjzjHz8QUoOKYkYzbbc7ZzzN2m61TiWD0t0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 107728)
LBbevY9tbX/IXhS/UFWfwyT3hZnREU7qsRBbLyvpNKEhfe+hZC5oin3eIKXcRDlX
gSys27zo0yA8NXrOHzmcMeEzlkVIrvdjKPlaXk6Li/mM0W9y6e65KzhQJhR4E095
4j2+1dPGgWyPbbRHYu50mAiWehDSJGwUwu9HMzPlAPZhP4GR9LfNE3Z73fU2qsPl
VcpV2I+h9Q0kzak5w5qdb/KQOhm02jsQ9dPtrKeVllh1cAmWNGWePnppUaur2AUU
uq+GKX74wdSdk4DgAQlHUd07KwMGeAGH0npLu+k/8iA+ENy0m5pLqc/0c0XWuTZ4
H9X1OcCDlP0C3K68Ou7fFylCyaaVeBaJf748JuVHHuej4u3H1y1MekFyRpTdnp+U
ARaZpSUOZAdQVCRl7G6E+Q+Ft2+uMWh/7wBlReARTpQiey+yN/XPex6EUH03q7L5
RP+du4s/Hi+ks2T5eGUMPdy20LTyavWEulePqaVjZxc/nVhzTp4OG702/2Q+29ym
XFUNTrVZ4XziSnLGuCBEYczXQl1mse5s86q9cUpy8ri6Rhy0fMV7hl+ynLu0hUo8
CsGCwRIIeE6QMkLtoygaRWWCcgjykdBejKwNLeq7AsHjfBL7r+y1i1UW2jbP8AOk
r0MFNxIRKmLpJT6FcwZTDXLmgnc1BZSPgmPOVPDDCMR1WpHjJ/6VdH/xjhv8W6oD
nzLmwbWwa9DMu8XIZIyxurgK+Ajrgenx26Yfxv/UaYKRwsgPxoqUmo6Eiv3LnOHe
3rWS6HlVWiYhvfN8JYaR7M0Srht7F6vJshWuQw3SsX5U9axjRa13nwELb01N4YRG
P2ouOqVFhqdpGtBo5fLE8DfM/S3ueqvEdnNOLXMEicvUXrQ6CD3dMw3zrNj0eqEc
Tj4+kNXITuRiyrCrh9wD+AzRJ6WWYfPPDthECNeY9BX+LpZikuLlgipv5iwy/OFh
cUcSKZT6vnXrPjElFzbj+jslHKD+77dX5hsr2jdzPUnK7z1ybkShJvfyrfd6/zwL
ffLmm6jgOeDrouGyJ0kQNy9WksOPPxhPUJGN9yRZ0/bIclcX7OJJe6qynUZSdSyv
JPiTYVyEU5dTFtKcl2LyfwTqJLMqbfsKOVc6sXYFG9xi4n5RcAog7iRyXcZQd7QA
J/eNRFoxKUFJVMn8kfEhaeX4OYASo7l2Tt7vbcrBq+6JLv6WOogld8deAT4qivff
LZPg8Av4hstt+40kUOIxgVSFDmgeWGSaDyLSfOuMJBoKh3s5TItlPnW5l3CB8s87
HpgzhxZY8tM6eSemZ2V7OBq20hwWQNN/LUg/IpHJZP2GmzU0YQCJtMQSS1kLMzZk
aQFYyWFDOxpa7hhSP6VHHZPphsaMrHj5T2m1zYyH2J8ar+Nyv6lkDjwT2B85SiWB
6Y+I6lzs6YnqwAuk50kvQNGnlsBXQjNWovQS20teZZNP3Z4DTQiu80boDz5vr0XC
S9vg6cgTVEDFyYci5tyEI3dBD4RHrUXYgT93aOfvmwbUpJWRvXz/u9KPztILsC5R
/StlUGSqgcbxBmXLlC8yw0L//RKl5bc9yuIUCj5GACExls1ozrUAhgko1pYGFxs/
HZkVzdnD7BYJaZ4+DmqQaLE2ss2mbgGxlFCYeDA5TMZ50CIjyGAisJCioNIt/RFX
I92ZxbRmy1qP10KltFPRxbp/yvcVEkEDE/jg3KpoSRN1MkyCmuEvoygM7jXGkb1W
h2eJFniGKjU1jigmwRw14hnVfF0HIvQjaMxq/uTrUOpDoJw9AGdpxBL7/LxqN3h7
UtJCfuuqAMuN/z+G2Nm016Pkl36xAyRLQ0//VSObKFQHJXkfWNal97/PE/i7RODv
/XxzHH/T8consgQdTYo6wLkLFYSaopxM+bDlJk5Wn5FMd/OhSe6fXKU7Rp0RGYUn
UYP4h4o2obmSVkwpDUVwD+kobIGSAoPY+AM+RsYlutg4fmU7AeimDRJLjAMrwmxt
3iTqKDO8BLMCeRfLvpIwQuH2H4zwJwQUAH6kLMylZqGPCuruJncV8LIgBhxZrFah
sHoOW1+hqsC7P+OxHfSLfY3hlPPAgouJSj6Shr5s+pZNjvDNwHoEmH6WSk5E6N6O
pYJWsTt/UVe7bBNKL8jE9vwh8QC8P2qC4cZgj2jFUAf1qwA9HD6oiM6FfRpQariB
+Is+UUTJWcnO9W6vSnPNTTtDH/4OX+HqdbrX00mplVIelJAPn1UPcdtFiAl5MhcX
fhqjiexquaEZUzssUfQYr9tidOAVJHF6sR4BZzxIO+kSQ+OTNBAhrBs++XdMoG4T
yi5YMCAjigRi7NuxxUl8IGRzB+P9e046SGwU9nXqKmE9rEJLUKZnLaiizJCxrO9k
/9GZgYGLwBWoRxOHg5M8GIQX/nt60UJIs/agf6yby6P6vVC/TVoVIVTe4P0Qzkzw
dIp5aMN8CTShiP//l9LutkbQQLD1jGHsyRxajk9LlA8L02NNgMTdEIGSX+aDcsXP
yQ1ShOvagBdHPqYQMUVRnfbLpFnMSfo/eLPt0o8+jnxwmdACJK7k5kBY4KXCOTMg
zvQTsDKqKM2/7Fl9rjffyi1zAPQQbGI3eXTiQcRY7dFdNTy0O7UabfOID5FvMc36
BfNhcIhlKTdXT0qbHA5fpZsb8VovdxINObowE3gihD6wEu5WLNrjT5ij3mVXCkqP
2pueOhehquvzNJ3WyBcTnn1fBD7a6ZqI7DLzWGXmTk99YFxH6LMB8qQ4fz6xmINI
DmK49OKNAL75cL7DIomH/fcngb+gR95y9mdsHPL2Jj5WADv1lpSest6hAPgUPtus
RYTej6W/hZHtNgkX7v+8owJY8zOiYyYGj/CyA9U42Ba4i9nT+GZ+XDnVcgr0QJ50
zi7DPrJRrP9sgV651p4bUvdXglJC4a7SkccHLW8UGnciidO/rXP5TatQScqrKCsO
/H0ULJ4WHOTHhIduVSdPOZBYZDVaclo3zoaWSgFDQ65++uO3CCTWyc7w5wbB8MTT
g/jla5lbUbAqYE3ALaZHRImz0uxBTYWuqVbbltO/NHJn2MMLWWAEIYpGPtxImWMl
/YHuiTFx0PMFV19u8MaWRIHmg6VW+KXTGAyQEgQ5jpbFpO11vTbuEvAWNWn62DEF
tUODeM6DlNIeiBkTR7mbW7wouZ93/AsEL3XCVV+p+NNn7j/FIbdLi3jQ1EsL7CnE
+8l4g6QhVFTqPCrxNvcXwmEA/mrSnZAC01+i83JjCGUtb+TVlWrUsFOwilPJDqS4
K2FCB/nHOswDBj863k8XMpmAiYLPGkuK70lsHoC/FgVjpuNc+ly+U5z1PaqAQ+kH
nZGsIqz73EEIZUdyoxF02sU99NBUFruvgb1EPsUQ+DYHaR3zV/D4Z/lBclyMdnFv
gc57gabrjlxSZU9Xcbfg5nbYKEj6/XAzxyWsDHnxLdcPuxAKbyi5SY9l3OZTP6pI
XUUWm/eaRU3hZOgnrogetLAsszvtwzhVWE23FEJhDH5vQyPdv95YWL56mlMxKTG2
uNjfzOdhNLw0mUZEwA49MrdbeJok6jkiJbkkAyIOOo3DqQn/DTvy1mE+PVP5ZmHJ
+JKBLQfdRS/4jhd1nEaIHS5P+8sCmDFtU3RqmIzea7pSKFokxZGrjz5iE4y7fn3G
A6e+yjY4gacWRr+lWVzhTggz3gGfoBM93UOAdIrzXAeaqzBLrecmcWo8Tbnvkj2M
EygCjBMJuNjcbA4n26MVsLImpUiZPcXrFsgnY7wcBWLBdeuJuS3U9n01tvmanbkW
tx8cpQ7ePkiTIFhXrENKTTCNXTO+MIbtwKYXKxbYYjf6fezDW6NuK2WBCS8oLXXu
V8whOrVMXS03S7TUinwwfa2ZRwhg1jINZA1qpnzrK6Zme57kqzzvzpeGAIW80cYB
JLkZ+l+zFPVQw0WsRHnZzVCDDiNSMF43DhCo5zgCeg1QnxudcBr7ERpwLhzeZ0r/
tZ8SVI4BdQOfMJZWpfgwiFqSsJmVHtyf1AfgXMsil4VLzaww8uZjXlCG5SLFsIEI
U03iFmwRohMTgJz8e5UxeCBlGCwdRqz2/kTDcY5CXexqGHaUvW+ZgDdGsE4W/Hyg
Gr4jb3IKbIG9RGtrtS9tUVqAfHKq2084eR7PRLpAUczUlvh1tQMeVHDggDInFUX+
LH9oPoUAa30CbdxBtcB4yn9lZ1ibSosD4Y2gMOhUTKqZ/JzVNhuhds1RTjyQSRHJ
gYsASSLyxU/eCnDnk3ADC3DFBYmHdBzrVVtra27rj8Lld+4NwXZXEz/+OYRHvJW9
ho18R6sgAOqLX/gZLLvpK9vZJGz1q/SIL0zX1iDabAcKVtJrZZutyh+OxeIJuii+
R1xBqUkZ9R/p+qXbEgwcS3Vg37CsoBwTaPWxrOVfMmoWj8hQ9Zhi2MHELY4TsXr5
pgk23gwxs3A7o+NJX0aPfbTYPWKYTKMuL83GssWUdyzzt48ZFEjE0QmKubMVko2b
tbmv70rg9nD0KJ7ugvJDnEGE8T+l7nMPVVUeKRaumLrQSNXbzAqj+KYOcmddR1tM
mG2yi5ZKYaEVe/5Q+wkULZrR/DCHIg0LFrHW2YJmQ7M8Ts+M62N1evNrlUzAWzOs
cIOqXWdSo4HTJDiS0lpsGS7xg4bXJTQ6Q3C233jYe6FEboZ7Oh3rr/6LyvCvy/kg
DdFZTqsD3JtA6NhV6TXos9QW5VWcisbfI0OWD99/RvAxOqHiVzUMPZ5V+7pah5X4
txz1KLxmhLvRc9aqqYv57xrhnQwJDoGo1XzZfiAuKkKus0YGDnOKqe+YUVyIVWbR
xcRB8fERKYnLZVc5YFq5mlWQYy9sZBJEmfIw6raSR7Lda1ud4+UuONQ7KAYVO7yX
86rhnspEQWDgyqauupHLGZsw93/Xn0TGKvX+37Me1aZ4ul2nXVHC/MFoX4mamuRX
qrjQdWnwDOIAoqirUY9ICivPUsmUM8CquW5K22Y9eOHAxr2k0uY+zo624YFUFyDl
SiZxbyt2b0ZuFMmKP+tPvshDbxts6lsgQNp/Kvv82ScIP2pL/NKBU9CDxcIpZ+xU
qGZ1lCFsPbfmznST83pWONCW68iuR9BAWymo670pER8KFpUL7tUh+MJ0hKz59tlF
FeGg2relME9wji+kEZeNeOyJYbxHgFOkx1puv56VVuagcn2ngVJkIgBtUOYYVzsO
Ew6JdC7d2wV0l9CinS1nMIRpRrslQuHPzClvxCrdHy45iqeyktYa9MKx618VlvOP
5bK33pN7hJMkct6nFOD5uUlN5XQGgP2Lpv+3dqERNvcNYuNNbAqBpmErFmL6VEMv
chDZstBYPdfqtlML1kIBVuhH/ehdIu3wLnFANit2L7438QNFjPLahEud2N18vYh9
EjTXuJgfaa4yuwZ3nRJ/ObSIJMCXUuX/V8Bo8GvS9b9clUnkiMmpA3XvDjhNHjiI
25BkrgXBhR3fwefaFGHd/QTXXFtQm7FWbUK1jRcpXeBCA8pPy46yHNe2l3Q6VnMK
tFH5I7ScjOcXLInuiXWtfLIiVqDS1OSB9VbrSKEUommc2+DReVIMH2MPIxdirdiI
S5e3dtnkH5bXbTaWVc6nCZZCvsgkDqGtOXfcZxPJbaaRnyFO5hB0T9SjnS8qVyvS
moz9sm8TmrdRB5bHHjxYy4XC3zzn+Y4HGdG8c2XXqYAei3BIeQu946DknbU4245h
l/w6jsbT/bxWScuchlqF5ZqHRCqHKt1OAvdI1luaa7GOUKRbM7P4iOlRlbz5bG1z
N9r4+X4I2212LLPl0wH+zCESH0fBh6h0cxTe9LM5gjy+wkN2Ij1rzT6qEe/dkDfJ
6soPSdqQYeG2LYLRbOB9+5Pz3vlgvby8lOAwenT29xul6daHyjxN5Dl4EiTpX4UR
GLh9jvRwNIzkELskKZZbzwFCJVNfvrfrWWvTzdrWzz70lO79uwfcZ34F7GXdHqxf
WRtPiAcvb359+xu1NfFjGTOXUTtP4Z5BuX9TipF+UqSWehdJUBJ/c1HMKP0l4t3z
8+lEKqD0BQyz0HM+4GOVR2MgKpLb+qOuB19MWlVZ0Uc5mrLxCiSiWLVcWDq/RuvD
Edr3WVKWBpd/6S8TMnirRRwqT1cUkaCzjc9yV16YcYeiF1LbutZExgeCUYfWkkHZ
uSbspbW8KVSZ+6ConGKIKvq9BKdBuclbX2Fon0REsgaLXKCbF2EVXR0+dyBkjD6M
gNwMJITjWJWYsRnUtEWBelvhuEt3Pa80MSo/NcV9tZk/ngaU2BQ4fnZUJiouh1Oj
OOBVLMipXJQdi4KwMkvvfLdWVQwuWvz0ptImVasqTNN3rAAZ+OVzYtb4SO5GMuLD
DYCYqpRe0q6K7keaKMFvHdZI9ujbVh9JPz6yOKv/7SWdLPteF5sjPoxuE99DyLGB
oysseUeFkCFgkvS6niy+JDCKgvwcJwtyw5My0lKgcxcEY6fR4GKIwmvXOaiYkUlh
5IFCqC7Ye6pehK2PPgzKjcUvt2YuutQbfvP4PXegGP7iCJsodA3K2AgGvAFWHPC9
lyRyPGrUVicr8EMbqwoz5ChD21uNBzP7l0lQy1px/UJAUIsdXXo4xfMkFQUpvhU7
W5QyjOPofCLyHcRi2hPd9pnxaLsjLwWn+GrdtS6F1ysHIq5Y6wJ8Wy6F848E5ZRY
mdMx6BiFDCS0c/3Q1EBSOFH/CBxoQ2HwPl1q563+kqexS5Y07/BA4bRxMulH4S9N
iV9a6LkUh/vXE8rGjxdpyg64YMNvenfbbSHmDQqf1fuo9nhgzKPlzATYrCORueFV
FAVRkoCGFPn3nnRw60mlYml4riDdlr9ulCqL/oX+XdQrKMtF2lLuxThHSj04FkdC
x0uy84sS53taKHv9y6ZhwTTeGDAvl/xBDRFV1Ve4JEWlLNlp3HFPb87vigY2l1O5
hEgNW0BZXsxDAXJvYL5b4gUuTpYKaa1Z0L8Siw04EZnoLXgX4hQKe/iTmG956zUl
BURgJ9nWHe36KDxRj33add/dkWeAilxxr3w1Put7UoToswupW7LTWmVvhL/3x434
YftFtpUcDPwTbmJaYHgX33WW72lV3nJSmsc/ToXDjrnsa2z4I3ouqrTInEjA87KD
EPqshJZF4Uy480t+++R0qmvM24XwPVPQktgnBIk1b/IttdqrxPWt5+g5GS5U3bUU
MGY/1sm3ra+h6dnqDDECgANzo/2W6X+otPHysV93Ll6DhqoydaU0aB5Sib2lNzJN
R4aY+I7KkGK3QWjlMHQHMDGmtQnGoC3xBPIjyYdCb8uxuW8dsSFqh23GtymsDYyB
TxyuVwqu2vj29hfkvtntxPZderPbCOXCGwv/gxbl/YCaWwe7f5UFH+v4jVOAPfo0
Mf2Q2Pm1zHBAAPjDS/imUJD1KOS0uAjZsUAN/k6s4S6w49rtjOFrlmlou3I2LUlj
KW0AMBFrjC1KTYbcnt/CFGjC7e2wOsxN9gdFHeIFNGSFucWuDR8eVC1YdVbNZMHO
5FYgPk17kOT3W/FF+ATYfOYp8KHcAuVmlkdQxXBbgu72ovbQs5B4ysOKTHuxnjF1
p/+9kJ7f6uSuyJ0cq/SmG0uka522dhQz653tM0ANaKMQLhLbcn/LoCPjBbfsFozE
PEI0smSNPlQKuYWtna26YQkYzAfsHZq6n2lm0Ah+kA1G0dKntSKPtEPCI5MmGMfm
pnTm4d+0GsCLGDE06Do8I5k1ymr/300AbPTLt1h4UpUf+Osaepv2gTDC9VSc3ew8
P7E45DCQ2ATaO4KbQu8yaVw0/e9XJf1/Zd6ZIeD9wbdX4UMJ8gpjH5masEkYA8lb
ex3G6OtoivWq7Aoa5Zhq99lP4BWppZ/c4cscX/TsHWY96NNEI6gsA+O0EJPc4JFk
LnimkkU8rijXrohjjsxksfWdH1jsDRWq0vZGjxS9dLD0ECXdn1fl+Tu29FjqboBB
z9j7iw1cj5/B4oA6p5Afh5MvXHKVxm9N18zenSdS9gEliZ4y8QZTb28btgUSMFcI
gBROsmCTdBSPWYFrutsRZv3pWfxlnNOOBzadYUvADQ2NUG/I9ZEoJAqPZfm17CWu
OqBF5GshuowAVmvILbz+RWUooUxNUaQSK5PKavKKSu/g3cii2Q+DTqXWTG9D7EDu
tqpgHamIJVm0oz98C42U7rXf1yh2/WmzGIS5OPivFtawqszsXnWZYWsKt3MsV7Rg
ai6D5VnAfPR3ok7u0LW/DPHwD+cN/ORKqN0THfaImZXALeSQavlm6amP+oFG4iYm
pvVLOHO029xcgq5UVnNkJRQHUjb0fUerb7EH3pPkYLH4QWQJkp7EiA4nYR0M9alQ
76u4DSjHID6IQdflToLIYqNfOhNMgOjY/1XjyYrlx+fN1QpVMgisBFfy6rHny0Nq
JY1WIbFVRIyqz/YdaZQA9uDrmGaEFEoh3oyN+v8vK7IigI28gME/EMu+/DhubdPG
B3LvsEzoBdcqLOpPtZij//431UhGbI7ReIwju3ZLROW+KeXjtQyu9fM5i73Jb5Ml
eq8qZjNVqucdfRFpwH7dy4SQklqCfqwJlv+Sx4Wd/jOoDnz52g+bMz4x4OHgsEwQ
9cx1spPoE8/3JSYYeDG0K31YNvjabnclzobBEvMKbwNTKSWyKOygNxOTXWmQ9VRf
GGPrRv0lu0Km6IzIUPXLTSAUBY4XC8y66rAT5I2YFvDHDmImF9ajIc8pQhRwjO41
mV93KrtMrpyp4y4azu1Jx5OOKZPlgeP7CDxl45SOGJKJnnaNtHH66mVb/EJVBYPW
8KXLTWvremEt2E/UVpB4r0u3GSGvBuAS14KOzQnhpIpJiWw1ue0+M8QzFixGQgmI
D0h8N1Hat/N7A/KoDhGZNWExZFImq00hoEvvN54a+n0urHSRqi6cmoApJa3K+SQr
0qZqYz6g7tgoWbr1q2tuqREfNTU+i+eVBfDJ7bUMt9CdEXpVBnVt2cKCkNK4nR2Z
8lY1A68x0T1w6diLPjXSn2nFiRnMipdTeUCF1/EUJIWpkWsk0uvxgX1gqTP12vGJ
WuhTHvFOPGQDR9ucwB27gSQB77SqFgYCsN2SsWiDQySTa58vi7SJ+1kiE5Q3ZaSI
HL7i0D4QVnyKPHfVDBGF+cV146iOkzLR6axUYr1XTZ+CexCzPIKjK/PGHLm1KF3L
NOkXpFcnx+DttEBXlJdlGz+mh4RnYRniTF5SgPrqGgtD+KfJWZgOuC1ATwgMeVVi
GZinoyEGGtxVEzQRC+zEJjvJh1mRbAcTCcAW52708zvFlPegOyZrgkh2JbdVnIA4
c9UDGruS3FP6TzZIAR5PK38f1fGwQubt8u6CWROlinnd9JHLFBkRDSSgauVjvD74
eiY6fyvvWanCWDeMV2YLuljhT1OhoF6XqohbOl5qD1xpgSPGwR0uOG/UkD/hSauo
JFlTKqu4ZXlAwND3Xht1u2Cr0RJq8t8IA6zG97QirCNzUi0aDSs64+oeKCbAT9Pv
/Wcpv0aN8ouUeT43mr0ZTaf6m/QQwacWQjBCvv4MM4M9ngf5qTUTMCaLhgvc+Ewq
lNIKTxSggqitEy0sakK8+zbcgMIkqafQxuP4iYmAiAYvMzSun16bbeXgCEYTFSwG
PIhS3l+8jr+G97NTFjd1Y/ZigfUYOrgqM+x9sk97LRiHsBW9f/LtmSMqQ4rcPme2
rT7bTxqlUh+yQ/I3BgUTBLehBQQkhuBNyCByxGXi3rs2DbE8w9bIcpN0y9J7Obh3
5b/DQzFhl+tmw8JzVI/Dkyhk0Gukl+BsqPc6TmzOR7br1lPvFO04Jgr7f/7s8Zwp
IdCKpy/cEQCETh+7T0DC28m9rGhYAtRVKJNvvIeyWwBpC5byV3EQy/wFut6Zhrzp
U59pWG+l/CgoZlNVGrn8NGeIo7eJH/AcZVl0pOqXyJjAt75xrEW8Gj0vjSGVtPv7
m7htDRogtgbFLBcuwiEUczKkHsnRcTFOBVAxObxojKb4s3noUC+ev4WOrrbBb8Nd
kmTf/UdXLMMN4seHSzvKy10BW+rAFTRZZklwyPUZpmDsGevPpoF+gG9wJbm1zNQB
CotVrd8BkByMRrKpR46NTs+2Csab/Px58J7LlTQylL/k4jF6v0nZfM/lCdu5zxhv
Hj5jyiWOxAkggmclMBC0wfEKbrTGnXpqcuFXBL2uI5dDjSsV5E0NqIQVdXKUYJmE
wx99ec95UIM/id9Tm83vb9WC+rBZczE7plUk8qeSdy5yN3trBWnkSw7Mmy6Kf3/W
yM7c8dmLVuhFiffAATE0UOSbPXDdpCvmlnx+g1tes6NkyW2k8tJEzS9XQ4j/7t05
39xyY4gYvIH7OcZb9ACCamv3ZkIzuV2oT1DXiMIgS2z+ZaOnuxtONVAOgYYld6gd
8FN17p3w/UOBiMkT4IZzvSQVv2WjPDkrNgzbiYKxDXK5Q39A+B38pLzQqG+aJYHW
gu3TML52th3iS9S0EMiZRwtgJB+Qmw/I57qiUZQ31okg9OARR9+IQ8UKlOyj7QdS
k4aZERTpaQo9EqLxsZZGsl2YvQccmDujK8dtZ5zIyuNM0hz3sOwuyNZqXwLNdPOZ
d39Kfz73H66Cdr+VLKoHXeKfEg3HE82/y3Qjy8/xd8jkOJ0D5gtwmC8dgPYTCzw1
bzmAcsovn6axJJmC6r1rTklTl3udj1RVBBAtivMJ/sjgdrACE+fs6nw7QzZG3XaW
UUNeiG/CmWyg0h+7K9OogpDA0SSzoOdrkW+Wkzsu9yP7BjNNnKwNCXu4NWWqAhI3
mmo3FuMc+oHaW4pfmunqIPpNc8MQI9EcauqghJDVWLTUkgwXJzlNqw49Lt5Wbvtp
RHWugjXUuQoTASVmiZYde9lcUQRFJ5KyqQcJuNBdATllOJ4WaRp7suXUqPcLhgL0
O1gImVN+UluiNHuTYPCWibpDXT8ddeKIOB5Dn8adu3Pvs0cUqH3To3M+b+t3fRnQ
GJdvp/u+0YNottPGblz7L1p9ztVKUpBTsrpEGBxED+x0JHhFqeFxi7xfUHrsWHeT
UQx4yhEWuje59V3O1+OCHRwdAQvDgj2dPMmSeU2cIhBunwEelKMy/q2BnVRRoK0x
I+M/RoPc4D59NSS+GjAbBu9f3jX8mEUz53JmW3dMxRdqSsSzqi916dg8ekgomz83
+GevHa+amTiEASIsOa8+N8f/ilywM4X3pmagj7EY4qMoYxtEgb7wBqg6dz57wmOA
vGifDQVVvccEuodCIbeY2lP3xju4x7iaPfuoazHBPzGShNdieDZlNocu9VuVcniM
dSenr2TO/Sj5au1kHI+rLtGziHd++uxaJt/W7SnV+s8tGxSyTvGj3MfZI6c16Y54
L9V2xZx/eOXBq588iXWc0ttnwUZld0eNUhIFJj+PXw6AuGgVq8cZqOowAEyxSvwY
U4faRkFilqjMXJYpPZFHynD5CDgjzgiz+lzJeGU899jHTP0FyauaWN6igiARR1Qo
BMLTFMRXASUZj6YltxJGfEsl1kQ7SgVXg0itm3ktfxwpRZWwXU7m7f/HBLotkA0z
srU+CBcP9ffxKxvNJy8xEgeeiD4FUqXjaFuB7LsflMmYh5BtoHVvb7KZgLI6Slte
QrHjuwVQpJQT7ooq9TzNhnyheQzGPw3M6dyyM8gNAXAt1JiyD4y3rKcUSoVqNxNj
lorrggO37lG9FanQ+gc/GfTHq/o5ezhMWde4aMR4sF9h0UJGrQ+EhFIOS9W0jH3K
PsH4Ta0hfNOAWp3Z20yhJD+nY7UeAENzvdNgiuaUiPDq3dImQDAeZtSzwEjiepZ5
h/jOcuYeodU65i9GV7CSM3PL8pEW0PyxjGVC8aCJbcKKItUv4Aufps1nk1qdQkme
H7U/5DVy26FdMwr9TcsX64ZLB2zq3wP75H+7uY1F3ZOQLqK/G1Ogf+a9jl9tuoKn
APHcBhwo4ezQmCowlm0T+xZFAzyUxllczt+kr+Jmp3+n7JnOtMqvizLoCY+6jVDJ
5a1zUOX//MAOMYPUhPbYUnMu022KE1T+22HAhNUtIxvnArU/+udgoEoPOxHbLCmN
uiXwmydFnoUlhDzkOluGtInMvtsHZZovbPxfz+9eDiun9ETmMSQfULwHQiWeaZ7g
InZkAEzdtlbIrsmdw2duq3lstWNhOBhWLzm0Ee34fVlFrf2LcV3vmUGOnEzTR5X2
qfeb5Dec15giCqfLBBpGoLJ3qXuuBclw36wL21u4zFVTwykZ06p5BZWtsXQuamER
89Oy0CDbL1jvodDfqkNnmBI7T9Oiv4mxzQiQRY9NRg6meJfVOevMtiaDHDcbYaZW
vtUYZDncSAT7ng+0apw0S5REcjiE0QTbbEQTsG01rtScqjEQYhFuZWI7vww/QUmd
VU3Trb9hRbKUUuXQIAyDkTokWgY2qnZd7G81BnewKmo3jNbWJgh9OPsBrU0qT8iT
GRQl4EIkndcl/Mr9occxvjvgdzlYsJFu3Ff7O2eXk1Zr57SfR9EFjArx9iQcj3KX
5x2m6Iy7f9lui1gZs7LZhO9ZGlxlKUIsbJCebO99F3QTSxxzI7BnZlav1lwNGixY
153cT6i8I0UuUnxsF3k/YuVjvkwUDOJ98tp7xVJC7sOlWFSbf1T8DUt14wEahC7H
V1zdRXdTdEIOrE5LVgT8MH3Y6VzZwfhnEvrmVzR7hVw0u6GtM44WKpCbG+axX2JQ
NvFRhQuN/j+IZUPgwT0N0ZQts8ZjwO3EkdOP7VOdY9HFJY5otlYLr/EA3ytJbEtS
l8WUi2W9be6HZab7Zp2zrAb+mKnV88ksWU/uGWxzrNUUEaUrnmGvzSGYchs5G/t4
R6QQ5iKw6ckjhIzig/VhhlTrdclKoWpuO9/Qwu3FOghS7I9fwtGD31LZyo1KEF7I
l4JfFhL+QZVd//VuyyXOlvdQI3GQ0iaKmtQwazZh4GbiKN90D+aFSp7wTRGreUd4
RD7GW15QCkMQYJ0AXl8Ps0WPu8e5XXjP2APx2MTiJ1t1DoKIpu/cy/OcIo8eXFlF
KTJ8BvtryGXvChHD/YTVftDrohPXJ2mJAA2kD/9Bu7LJ7T4CwALZ9sV0DjJsJIXK
Ic8oQhzgxSDazea6v0CrZx0FHot5SBrKuLPBk0iiHNZVlvx48S2l4n5AL7oYcCMP
87bo6Coz+vWMYZSVQGyoRuTjeuDFbRRunZwYctGB111odetUpnRjJ3U2hhCIMDCD
uj0sK1TM29vHbEWI4JI62vb9Gg87bnbxQvnIIaIqSWjfCFkrezzLnBq6HK45Jsqu
RoKmllb8hztQrvn43u62rS5FPIVRnl90oQNpm7CBWyDl63rS4QtKShmYQBOY4M64
CV3MLOkpBNh8i8HUD8ZDF6l+m89chJ3Ecz5vihId9miqWI21II2sRp1LW3PyvIwp
fEIt/hLo5Df1/UAkoafXIjS8KCiNXO882Pa5RaC4Ud06LDzfbwjLKNs/+EUoH9QP
tX+uStkRZqxcAMi2OFPKXDATNOlByk37A0ad+HnRYE1j9mvTIYPS2rvMs/Tm0MKn
WMVGmQvEhbJw9AGc3C0tPA3hqYcWPW1i9lpHW/t4gcpUvyfUWht3Y7e7IkWccdlY
gk+QslqK75GGirI6tp0xVT2owyO9QtZAQ6I2pftZYEECJdih1N8Q92nHlIUu3ODt
iZnoiNFNgRyfKoM3fJZa7tqy30vJnIn6avFFIUL0IZVDeB7Qsd6HuQJkLcv/LpRS
HNfgq9Ql8zbSGdbk/R2go57+tdfTTV4SaIBnpIpC8SmWnwNZxYAYCprkKQlobSYf
W8KGWeUd/y/Y2HoTUyBuqQqZUh9l1MmM2ifYSJM4a6S8wLDwQ4MMZENL+VZ+wVwv
m04B+M6hJ8ySqbVSaES1K18RHj/CKNADIy+yvYeaWsnqB+uCScYUmPq+awHqm57p
iuGUfOsDpFjPwSUhwgOPBVa9BK+d8nayKXDWxjsbCoQuL4R97ZtMRYbtW6y3VQNh
b57chWnk3yUDf5uOmqsFMjzUyuBjm12FAGYH50Lv2eeS/XFwc8K1pMLRxFqkYKNR
rNLayOV2iQSqHk84uGWhohq5b9ZU++ZEDMoaL7otLu+uoMAyO1KDo01vocnsq0rw
f01QHvGwRKWyWlc7Yc3a2gwwIieEz9AAKHslXTROPrzKEJA2AvcVQ4zVDsTPuVZw
HndmwskqPEEfS+XW7FRdEYCwcTjVDDByPRqH/cfdPiKF37u+Jxtnw4fK9Yih4ZLk
/iq5A0Be7aojLoxUcq7GflRfHnvQHr+zCl4hJnd3s17OVB6wDmOR9xVIQgGvGbPi
eWuKnIxptOu5iIaZQnacVvT4ELdoKVll2p11g1ikjxVbxMVL6w0kqIpzn9sLkF5C
kKn0rnXCcaxqjH3LTAaFlYqjHuwOWjJTL/+5xxDacUjDeu9sUGQkToAV6gt0/a0k
ACPh5fWsVFCMpte+daF141yO3WKChaGF4ClPfhK7HVCZQ9dsF8g+ohgbZhNvwviY
2TsxJso1M808zZ09oeuzgGZEgdxDO7+Xljm4PH0/Yi/RHeiM6KcNl79ZQ7G/i3R6
YByFy5rN5Z2NPz+ZIrx5PFeRSA1DxFAr0w/h/eBBgNnzei9O6+NuRPRkYxanWOUJ
jT3ZX/WLorWlUuCbrFbnoLLMdDn6eOyFEWy0EGo6Q8pghuJXvi1ZiAVr9D8sHJOt
1qj1zEvvSzQTLWmma8+nSYqufC44Av6ByaCW5nRfRa9qMHEW2CzB1NVkxST3G3tn
PnKDy0Fv5ACEswda9FC6mdNCgK6UJCg7MwGwKnOfiwwvC0T+WwkGoGmvTKRbQQlR
OcG9db4P5fWLl8YPe+5kMuEe+bqFFb7XyGKqaGi3VhEUbsKM7K45AZ8IyxRdzJgQ
Hh5F9P5QRNeqkSU1sVXRIU9CUA6wwBmFSQ9n+ImLa8SJe5umer9J8pfJtmZrRXPj
zzckUki2fB6DRnyTM9SRnE0DcE/uGHz0JIjezvnrGCb4f+YJgIeYKoiq1yhHhwdw
00NR+M12LoKYzfbyWzhxujZpLh2vQtsi9JEW4Zrkk5rz7YF4qJ9hDCPx3Y7gDgfV
Gbyeudli0Z6u+WAZGwuBIaHvBWjTs04QZlCbUz1gi/T/eKIdBROip4bopZEgBGtE
M3W8Zo+rNjK2+pR0UKEFqkE9AasLOp0xHCImWffq6Ma3Os7cGlx4xyNzfQz2JmUU
Hx3cRgitBJgPP9/ZyyurCU88h+ftDcnN/IOFZSDVDx+WGOgyYkthZLLOt6pTggfl
0FUL7YcKfWQh8Jf2Lmt7+l2t5pllfC+tog1Xi4eNYeTFXO7RXaIObVj1VTHa5tNl
/t1AWFlXlJUxBt4IrOSxzIMqAAXyGSZ0e1OAcUrZiAvWy0LOPFffOpF41Ro4DJul
7BVirbtsFvZFJsb828mfcDRJogvbJKD/LU+QYaZYJ5vN4i9iMyeQSuHLbvm0Fit7
S5eIc9/QUvY9NdkWohITxzIlnCgBO+xBOECGKJk2IOjQAsSUG/lFVidWAADm5fv4
y7wTPfnuYhIpVSD/Qo3EL0uEJ/AgH4DenuPWsdx7wjxZjPwToVue3ULepD9j3hGl
Q+ZGb1nWGwANTTZkl+i3UGmKvmlu5/EVUsMgy01h5MQ27CNb8BoAosShtkSSk4Se
aV+dwVJrC2H4IAmjxeTDQkQXzW8MNpZEeIYsBksCXvtbgBNoS5VS/gwKuAK/q/Vq
Pu7UiYaCCPrMsAjM/2x8Qp4hvNl3pj6CBKn81TU9uzcLVwoXjFMnA7BKB/98AzKE
dXTPvbEqYjrPQ0UlywuNAoYqQeVV6dF8F3ZZfC7Wocu//Z1793Wq25NvEhA+FCJI
HPa424kD0mktidT10UN8sxZumrbpJ0ZdmpUqy0Q8ITzfEkXfzfj8S0tjs/HlWF4x
u52VHtgaMVaf8tjCpg9zypYgD0/mHACRVKHPxmJKnf9omZRHqRAwNSb+4nJVWHd8
lTIOlGwWvSBm9bkIKUp6PvugaZcCJ4/UeMAQzA/zWgQCyHm+QIgyqTmfKvgl2eLZ
wJlx1VD2iRvAittq1xZb+2pWJd2+6jqOrxekjK/A/eB6SxUntBFYiJy86z6wZBgA
UA/ufcmD+a1oZOqdV59RoM3WCp6tc5f8tAWbz2lBEwaxKpPBN8ylAZv1pPyMr8Gp
7UKu34xgLArj6cHLKIsGH4QkKNgPoyoS/PX82N4DKNdktD9lQ3KVwmte7ilZUho7
nhKIfSee+i//cIFjcAtuM9J5fHZL+yO+dcK7l2SxOrxzrWRJ7MjsFv0hEOzL8j8+
uxsFoJkJwFuIwRoliJ3IiTMmxZJF9qmqKlFAvau6GQOkJ1CBZwU+gY2eJ4gZA9RJ
ICdho4wH0g+glTZOg9XS/mf7DPe17qIyZSWm953UxQQLX2uegZ4EIia0cJa4WUSJ
KgO8FUnxFQOYP68iYWOE5cUn5QxltKCTIPCn+Vf2+7bKY7IACBcSHTGIJfjnaS5/
Kn/7CscF6Ch5bb3XHcxjlkcDdz9UUmR2eQO+9OUjwFSpygh9To3EC2wHpps5AAD6
EvrZ37Q/Te+OB8O2SLvu4r8+U+Ce0kQgiuwpV85P62JleYz5nYXcVBXVz1eRsk3I
e2xYQkHFyHRTUN9wLlWme28gxpvLBDsYnqKTFHAPNPLSSAhkQ5eokaa+I3ZY41Px
l14Tqmt2821jeIqA6s8/cBOyzCsPjU6KyTtyTyfVahVwDE2w3M73akIMkzZTWZ/a
uwKO8I+9L0It/bhw61tbor09iU9hagWyclvMWFb6wyFZL13761n+v6V4w8pvuaNh
/DA3vOZfuH5VeWHSMS8yMfkIF7Ilr+MsQDchwNx4xNYZATp4NYxDX9Hnmk9GjKh6
/vqKieUD8lluT5IyU50YFxpzUXISx4XYqInBmUYZ6581vE3s8XX6MbDE5R0ghIal
XZsmmlfCFjZxYM8j+DBK3r2rwoI8yae/7gQYCDyyBviK5nVoa9g7emLXbXfvXs9m
VUoiaZ/4Ez3CwbRvimX1OIi6hLRv+khadHyZjb3FHIJc4+MjCiJiQz15DZnX9Hdk
WeqpQ2i0wDanMjZ/mrygORw2sxY7L9dns58T+AdcvzwT0Oct0wVqbdybQkuTLnfe
wFZhLwJa649+05Z4WMBGxPiB/9l1uJZIFKxZku54uJMYTv9J2NhJ0BLhsWf/zr2c
sedYMkii951goE2ml4DQllcYIkG/uJBR0LDTTEvgndwGQQ8VHG7Qloo9FP9oYVym
ooanCkD/zaN9WnANJaSH8JvvcWtzu1AJpJ0pQv5zK4T+Iu4jnBmFn2QYKwClXnKM
KI3nLE1x8ykVlXbR84Dm8LS6bBzIOD0m33YesJzIqdmMyN+6vLx59o9wbozs95BW
ugz049bWbA7YEye3124mONACGB+DmTCUlll6fIuYmqyjDo1VkbNS2MERGt/ARp4w
mxvDKH0U6re55eyL52ahUfLckpOvcFYgpxAQadDNTraXKaxL+GMOVE4PkOyFLUCC
63xrlPapO4G+AunL7FQC1yNMRXtniC9O/FPv/rRwwLVP7glzLFwF7n1Pza6RND5y
YjP5LMQhdP56mucs7q6VWKN2BqX0PsmU9u6IMaNc19JPLSAa5+qopFvDIngcMyv0
osTvqd9j9D7RRMVg125CwH1apivCV4Yo48mvv8JZ/gTLeIsrNh+tiJNKvFdPrjFQ
0xsNuREW3qYpdS1Vdm+UjtuVmqPiubd/hAXDV/Nv579aur4g2xP0UCiOCvK8QfUh
lQrLRXN6PjJ0IgHUwaulLpNiAFuCkcl3SnUW5XHSETmNYTDCOtabSqVRSnhILtvo
yMVdrGRAbByfEuw1tZ1MQwyl+F1pDhS7YJqT36Sdpe9AQGQKO16JCEsnFJrxaQjX
BMtORftjdswLMgdCmEbpcuGdOP+jYYK3GXvaBjVffPidgGpytFj0dg9ZnJJZD6RC
wLyWpxNkEi4Hxu/nctGx2Y7AEy9vLX0C6jcViQeXDfjzWvPaQ7T54mb92tBUs0oh
zWNm2U27Lm3M2GwTJgKXmN/vrru7CNnJbH+YHPNoRSFpGbX91ZKtlbdgNfAAdLWd
o9Oa+fZXxxxORbGna3NwWoa3R85246ZwUNTA6JV73wdLMcMuz+exohH+fPLO5fY2
MA+/gqoUsbSIgx7FTcmcUbjIpkCJ0SVOHv8CtsDykM4FcDQhmDQ7ZsXzINIJt7Pd
tAHzit7q+BK9H+hHeBtcz3Ki8vjpArRL/pR7k6EIWTOpEr1XJUWscTmA+PZxNxlR
+LWhHYupdW0eXEpdyZa+XwFhqnJvK0BG73kb1msc6j6qHWYeY4q0mXQD/wrN5gRh
48NyhoPtwsKBVByFQdFWm5Fp8wgAU4GMWglkOiL+JRo4qDDFQeQ3SqRaW433TA2C
Pef7o7TahmRFC8qdQuQ3aToJqsGRrGLhfa4DeNiiUbOeZvOff6k/ktyQYSqrJxRN
D0/Ym3nrwegnklem7T1SwH72kSDT6G4Y9SLwb4SWZIdkrxQRPzyymsTXhUdD8yEc
jSiI4WRYsKXalC1tYlzC8Ze6t0s8WSsO+EbIUY/zHRrVlcwTYhlLGrt/Pn4M4bTt
QxBgwbPNLSz7H+FlwEI6i8neXKPXJexjfQy9FzRwACYgApPoL7XbEK9g9zjvEGC7
S6WiBjzoaGb5nQKfGGK2CVciVjWjcr5YQHDnN3Dni0saOWbRM3qBXnbLx3NFUzzA
dliAMLNTr1BS5AugDV/rkJCPpNZ+7hSFHE/WB72f5NjTTBDMi5mu26nA2i99oOve
VAnaCa2pwdhWxvl7AUNPKtXUme+2eveoj6Tj7sO/ZqcZ5Y4Yj8C5hlKu3dQ/055z
CNu2OIA55uMQIW0kQL6jwzH2jMlrG12ft/HmtSYBnP0kqlEAp8GYIlqT18hnLGwb
1eSeEVwanUZW7BBBqZc2wpVjU/37fIVkD4oP/5XrRlFqhD0HB4/3JkP7zOmyOd6y
faIY/Q4xOWwydtr6//kpahHmFkIzejPSDZAqPlcd0kYdCQHQ7wmGrlLlUr8xirhf
6mCl5SXFN/Co/ZG4qN4YrM3il6yPmBJBbK7jzWc8YsEVV204zbRVkwgLFfAxtkXi
0wCA8f7Ckk3TLPXq6q9KIhIvvshcx8PdcQ1yg67rNZPe6b+X+wMnaZ/pxH2bCCbi
wgfomywSpOuQt82pOUtcGF1dTvjllPS5YmBalTCVuoMLSFrJ0iIm6w0+6Y3phRLN
K4YC69BIv4v1hHfj+YmihpIbjF5U3ksRMzB0SDluDR/iEz3qt+hg9DBcrri4g9MA
g6rPcpD3RMq4oM/b33zJD3AB3IQ8Z6IyJDvQsxIVdeK+V5XhSt5tYYJGfvfTup1F
fS9k6MCOfPnB3W9VQhTCr3+txCEr9qh7zYOkrMhJ2XnK33TuNbFGDy7Z57hDmFcP
m8UEKfc7IycwRbDREfZ8avJK1IMvNVxn5P+dgzZhwyTQGgC5fXW87WfvGkCioZP1
k5fb+GgyfOlCgjxNLpZtyTODmbcHO1MorEt2jY3e3qUBClaI3a1c48NnpwNHhg71
li8MzBaBjqDVwcLaJLaRXB3EanRjjhRWmm5DwAyzweW0gteuvJK18/ZqPW9wnY/P
c91JpP3jeatX0Y7CwxhMPjLRdx7TgwW11hYJmdVhxhhpoyVcTmQn3WeHjk/fu/yP
pcRNwG4NNyLnfFiydcJFDkoeW+otLPqeSkCGxI+Aa05qeQsji8+ufyHfO/A1wq5P
jORLnZJI3qUkFSzHoYyLEjwcjJZ7HHPqA9bHUop4HTh3YklGackYjNIsLC5a6gnq
qQvSRHcQqMc73dBdJZ7NC2F29Ve51XkLeRFmgSNxcLU8jI6rQmbfCg2BQGYYc4t9
p7mTULkrcfJ4WZuz/oX0Rw/k2m6Qo/Xv/vIoFbSIrCDx7QARn1D5QVaGHayFrGJH
iswww7/IDsWX5XPiMLy/wpVf9WgZ9MsF2hCeVSLYGL6Nq0BdLaGg6JO01R69ikk/
e72h0UlQ/iMZ1wfNknbc3f5FcoqHQhFXRIkr2k17HxgJGfrRmeJMy5vSZ50KjuDQ
WjhrW38EqQI7gI+TQTIXx/yZEpm1BStww+WJ6kL6sR6pqJGs3IPWVf5npVJI8YEK
W0OXhqkBauM8WDgu5onzFA2y2ULVknng+WvzFX/31ISq79mYGcN70MwwC3814mUE
PQZAN03aAlImDrzSw6kS88He9afLlF8zcQ6ErGWjTbfl5e8haZqQSxQP2CvTcn5t
52fx82CL35ack2wvnpQ0NM4+2+olJbAzSYMbTOSlzS9K1Ko4deLwg4uuCCtgnfgj
Xgv7LEZYrpeUkIyKqfWMOU4E4EG+GiFPuQAMTCXyGLFmkYwHHTHri2EsxTButLi1
j47dW8QucXjnmWZl5wAkw/IAbHQ0k3y3N0vy2l8qvRhqq19uycxC6k0dhJmYtrf8
FpbBKe898VXeZaSQhQwMioY6ulWBaJJO9CJQDhGPkkCB6a5xtDacuR+u8bvP0OIg
t1DGYW89nsInhGZ+FPQPr8MrkwbSBAGlZT18vGqG7gXnTgg1eOxKpK6x9tvbQYVf
NrA8LKO02fVxg99e9GbYko74gfM4VuDeGrcWLEuEFW5FEZ/7vusL6kXnGk/OyjXn
aS08s8+v5BaYaXts3Gggi1a3Ihtzqqmfwn3mqkgU8yGrTOT/4Fy/IYTVpP+b/4Ax
Te/kaV5StZ8zB5kqJq0wuqtqTgKoE8s45QpTZt4YKT6F0KPHFvfRV41XHP5pzjc3
jJ7GPFY58TOeyqjvFSwHr1SOrpGQ/DrQ2nTgTj3Swg2N66yO/tr2ISZn/In5abCk
JK0HBtdKuWL6aKk5vxkOijurGlKmRcwSbYA1LYoPsRSZK3SG7/6QlI32wso82TOW
LMp8AWLNknA1TPgnfbxdPwUpwJGX/gjSsqHrNmpbuBLu/RBoM/ax6FdXC189wudl
U7/LHv4XLuZ3p6a6ZHJdv8R+PB26hfVFk+buj+anqrinrtg/NIbg+umPfbl70dVa
twss+TMoGUYNNtlUaA994F+uE9M3DTvl3ljrlVPIRl0Hwbg1D2OyQTaA1ziUVpNQ
kxuT8Lu7kk1Wtkv7II4GPHvxjSVF0B7Z4z0djnwx2wBGbHbrQdrnFpMZllQbIwbO
A4pIAI1e0Yp+3AvVIcwrd5sTrmoEHQHjvJ+gOfpc0U3Cg+L+PAA4kvOPGSChewbv
JCRy2W+uGG6QjNGxxQWiFm1W5mFQjtB5KrfnAOUmKovh/J8jE1wzI1fulDFDnD/f
Iec4RErMs2DNDc89RmSQ8d/bG6LWFK8CUk97BerCsZU3LOS9uV4uEnIiRQGLroAs
IEBTcP4CcXjtQ9sMGKvfQkqSuktAGrta300oi3jEG4FIz8DzuZTQv4l1TgETcqA+
T6L2mMKCumtNQPlx860dEUO5bwhIHKKatzXiCOJtd03t1leqWN3QP+gfks4IjJk5
TMA0FwRam0vh+VAj9YHTCDxOfodipUMdG0XAsm5XLRwDyCFYtlx9x34p3ByQPJ3l
6QMiNKZ4/VqT46NgMGAlHAoa4IzH5q8Lh1k7jctVt1gBBGPDuRqgQqabBNOAnMD8
JrP9Xb/cbeh083fT+HrtdsXyZpW5krCLTK3qQVWf4RWcBM71EKwblueE7nSoN6YW
PcvfH34YbYPldRVc0CtNguQCfZUqNE9Cplp4j3q77ms8msjoRvFCYJiPzqp4yVj3
e9RlvxyghZGNuJRxhXbQ0FVUPtpouOM2F6qHHsrlGOX9Q89s7FGgUOFwBNyYUPo7
tft76iAj+MsERZylleGSMJL1LoF1WxjfQQbXD2PUg4XFqAOzXzuJpfK2COcosaRU
gfYnQ4QAbaAycB3eB+qW4577PCG7pD8N0vm2T2uG3qt5oRhv17VZBVH8YkO89ZqZ
hzMJt32OgRnUBM8LF5MZU4wDjIuPH40vWZPmej0EwnHjgAvgO5LAWo+30R6W/Vbc
CJm2uRC2AAY0eEmx4ENg55/W2XEDjVsaupCndefqDgjdBOOIvJ7yQaUnjGm3EXSt
qqma3Al1wE7E8AWXUUo3eDLPx7zWzwY+1NSgkl7ief/zCT/MN/6maUpjMUHyEgmK
lY4/zYpRuQmEhPLLqKDL82ql3TNbsGe6gARU7u0Id+2gZepzn/o2vNjM+JESzNcj
RJ0WNhv2oYDs++8qA+qS8lav74Z19MwdJVpN2wS7BGbRmgp395N0qp3Iy2BHRkcl
Wg1lNHrMfaV0TE+CJxOkxM3KIOMXzYuMGVrDCaKLvaWRpY0kutP8vKHE2O8Cbe+r
9gGlmb47fLd/ZdBMIzKfNKEeCKqA4N2TLjhi/chWj7PnE5hHF8iJ9Omq872lbl9Y
bEDOGtAS8X/DldXJwhBxCVlzsxr8HEY2qQaWCVg1pPXh2c/gJ2JFmQSAMpvA6wo5
p3M35C7Q0XQl8e2HQmJWFeV8cScrghC4DwFlTCfbsxvjvmke4KoC4LTCAVrIOqSX
R0iZGwmmCQdfj9yrc/Dyylei3rThZlP10t5iInH8pJpxYQsvfnIQqtFELBLBPI/w
RQ2m0aEt0DC8oDXd9UZFmOrzPUM0L4wuzczAL7xLwpzgAoEekeIWlftYbWmq5Juu
RNpWRhsUKMklhB6246eYORe3JajPobsh2b1ABZQIeZ81a/i5Nezsvc+t/nJ0c97k
G8aRQ/v6MpbeZC+xyhkiRloyRTE07+NdlXOYtyKZjwy4KiRqUWxIsuBYlxgE89ef
iLFFB6GRIE0HbuBYTPr+tngX8BDOb88XKO/pQaop8wST/B2bdvyULN2Fm4ufZ18u
Fl3KiZ7o99c2jZFNHI4LpPnozaV5hH750+5ma5i9KQsNOpN9VVAwWY6Mh2jqoUZO
EJT3K7iRTMz6sYbRXSOOYmMe7PbXe4iKY4Tr5Hb5tiW71PV4giZfIyHvc+k/LmCu
mseBxmfpabbcjBieuHlF/wjWgjNzF8/Ui4MLWceKTUOqMRhgpNCQ+f3xQ9bKyltR
BdrLRPMTHUhDsr642mMNAHVOQz7XCEyurZ8HvuNYFGM89+ZeS0w5G1Imayo7w9to
4Ho4PVsQJVugqdLfAeTZhdBcVhUI0NEtSv4cfv38xR6t9eArx2gBjgiHTfI/farT
75ECaJtbGW8mnxPi3BTnPghNo38RvxUllm8qqrQA2aPO5YgLwnD4+JE6JnEAYjFw
zen8b1e1jGgdFQLdvth0ABF03YFhU1K4nHsTITwscFZIZhymbO74mQ+ao+RxiSGz
yF77tPh9BnSmPkFH23StYb7TUc93V76SifcHN1C6mshFQ/aEntXCuDp92sImSfuY
sjDO90kSzjdUB91azIk7LaOorbOs94HkjUDE3/NMQ0uHtLu68PY8NoySBmQN19qu
2DRufjalY3nmHZP03dAiL+EvIWtGzVOQqdWC7eYBfqByu3U9aZI2VGSnWD85cD+c
FpeNHc/KgbX0HOtk/qIEqHYdXKHckRoXz9CG979/BgGVynRKE9M7NxxhcsSRb6od
Ydpm8mgXrMv9DHrzVlmhfOjs+57gnOnKa6WmENn0ILzZUIasVafwNMlMcQb0fZW7
UjSnhjgjqRb3FBNKpIp6DPMNgfwOsyF530jkL9AfI+o2JguQZlLFeip/1j6GdZM8
GHEs64sUg6YenQcjz8z4hgBDJ/jWijFRKW15LARKb9tx9gYm7ax3ELCXDboPOf2F
hoyhmj3OGI6Np2Jtj7ORXGZlVyIOOxILCGd4gY9XadiHdmSxbzHAcJve0aF4Fafg
tzEpKiZE7hM0lSlq13f4PL/Rsk6jLTUgbkbW1LKJ1WXIagfJOWJl3ie2cj8OvSw4
djHYaV6J/Bh6L06fcjS6IOJGFnZ1uXPrW0EwhbnVV6dK6YPFxZlrka3M2T2zGvgu
2CMVmlD4nHS3TGZPWgrAQrsEfNbzsje78yd67Lu5qo6n3gP70fqshY2N9nMUVGBR
vMveacK6wm2GeIgA93wYefObch1VwUKX9xQXeK/YDU8pZgkzX5cn3tZ3mvSliWVf
sWu1n+DQwEn6l3Hq3lXNEfbdZZFl9O43+gUuByuTY0EVTuTrlKpI+ongHvI0z+gz
m+DTQZ8v8anDZYbHw94mZJF0efJGS5duyaA1wqTys3Lel4unpwN+3fgC9cQDLJ3v
GtObPKl4RnR6H/96qWGO6PMrXZLrIKN9d9DjhF0GxBSfGF6doUG9yqTp8M4Izujf
zWoviz9aRDm2pwgvgNEw/Cywl4IIHszi49d4h/dCfSFzC76CTRKUoKxi1MmK4sAp
rYY2X3qF592su1vACLEoj89ONcaKk+VQukvLjWTtowCG+bMYjXBNhV/a98R+ox3M
L9xUahIlWzA01nH/fQpPgKGQM3cma94ZP/IowDpw2CKSV9C8pi3sc5DOnroy8Ks+
2iEgKch8wzsfpgY/H3qu5npB/kZOGL9t9qO0Ka77+0+1NoS/63ylUwDgS+cvl1bI
+rHOaUeHNa8mvgtHWrVEZvjUc0kmWp4L13NxP+CKS1RcXuibX/8izRdu7JsHGI3l
Mkdso6eibuwv3YwR9kyQ35jtSaSE+EmdYB4lnNasy8AD8u9VZ1/JpQ5uyTK0isUB
ZUYpbxcUIz/LUi+eSFJY7yKSxWxOXCGzWlFP7yoOxK4nYl/nWpt8rNE/qOHkhaps
n/DBaY98iUhpcenuSpcGFDspPEadLFu7+X5jst12W18+mo4yGsTs9NR5JeexYWjB
8dD2h3unRvV+bxgy87lHnVoob93QTADZuZg/RyJV7g6xfv+Ek/u8ZKOr477paH/9
9EcCPhFDsSLyZw4CmJ4TjNXiKQ1ZYwkP7V38N0LgLwle5HnjmhPAL3WR+m686VR+
xxvTBz38i8y4RbWaJQDgskrNF4CiDrB6wiLLxA04l2RqGuiQbW46Kcmno15tRB2E
T/4vlOXKZggCMRr+ySUrU3kMkfImvJrbFgTyEJo9CPLj7zbVBv0I5V2pRlTxhWBc
9i8NHB01s8iFBz3f5GFuUZZgBdFpEXUBKdpKFwo+D7tRfsFMFvq47bMl6zAY9i3+
cCYhXAJZ6VgLzW3cxMC+JNQDfX1EnotRcYb7G8sxESz8wvqghGZmjIAZFNRhbmf9
em26DLXnLCC9fibQBpMzoDvaMsX1TzTuckXlSVVsMLpErYQ2FZzj41row9ZiEzCB
uyg1uz+rsnJ6CI1mm3kd3DOOM3eP73WRETemPTPwCfsoIkCpp4yxo5IX93TJeaMT
n23IEeIi/ApN340i4JUk+t16LA9kvKcqYRMbHzTPWs/ugYwoqhZxOAskEcOgeBIT
AYP1ycVbps7lWROcmeqU00aU459vDcLhfDKfixH4PDH34fq3E6DkAM++OI7GQuyv
YdarEjI59RYCD2EEcRXBxwHcTzgZLiKT7/L0V8GFmkL1dALvvXNYtFIYH/bBLRMX
CHp/aUOzi11ExNoBHBQS8OkGdvtl4W8USoxx0TDaKmOnPZh7lbrnNJCgVOoMpVSb
xxuZ0TtZSg3i1nP3jCMQUpGmn86oTiFoBBPDW1sIr1g110flmP9nsatYmr2cHnTD
eS0UvLl+A1PK7/Eqm3s3YGwwoXjbwWtSuIiwEbmOZV462ZDXHQE0fBSbNBKdjPRV
J7g0RupmdftIRamw9ViJ9/mfCjffAYMl/ym53fywqbpEgKwXnNhrHI62sKtD1XxU
WbI7n6/1bbLThRtbEDwPQP4jVcw4AmH0QBeKJyccDt52XFaFOt2zz8vwFqXG/yxj
lEJW/YBuZGzthEHC8oi8kiw8Zo9EE+QSxzItcKBg18aOp5oBBe0aU23vbpQ7iXPP
S3yWZj2+jdCiH81pgQrAoFH1/edzjA5xu+vvob0GVFPbeAh9/sjHe1R/LgNNKu8L
doD/NKst22vxYhwhBl6e1WRdoMVXb9zz9ZnHmz9SdJk1lP1pRQMbq6iOssQB/1Gt
b7pBoS7XmovJd6lA0uog2iZVRkM5TvogDR/GgfkEGXFQUCEqusRa/fg756TPo7si
ALMsJh5X9Pe16CiE21XQjopRPenB3oRNXAqq5ZAhKAPjtFx114fqi6V0fCkrwR36
Wybw4SAoALwzoSNVQzglsnVCEVTsFTwn7HFDxpKmR3A0Hlheinl59qUEKvCRdc+m
zt+3tZJoGM0Qw4zVUD03+cnEI+h8kkkOfxs5StXX9GlMC7hsm1p4mN7PBFJz5VbC
7hFH2ToYNCyNH+X1Tq92zU9acgX1EoPcOikPBXmKZ4GluQc8D3e8is001I5jnAy0
Uub3lQfOHRNTOB0fPfDPkIO4Cax8GOI+KI+cPygEudRvNAi/VZhg8wJuvpeRHlxF
o+/58SwuOAQ6sDcZ1M4Z1r6vUgEl/KC0XTAbHvJx0LiDCJ88OYdpI2fBUnBFMkjt
WgUVd9WMcN+WHPL1vNKtej87QrlojHlKB1XDWa59ytQSk6majtyZ7iedfmrGAe/3
3EiQS8rsCtCmWOqNTpd3MlB3+kpTFoOE1lN2XbnjYr3VeVFqEuGXVALx95WY4JTc
XibuU9kMaCLZKXeD9vVkiDqrG7GQgxjCtAtFeLLnU7BDYLa+HAVJfbP3m0NF8owO
mqlYBVz/XFBckHpHZ84CXL6ti/Um9dHZ8jr2QoMzpdaPlsU8Ome6BVX2lqsONXWa
RJZ+e45v2ETeez8Q+YDAR0m4H75OItzI6Ouk+7xu1BaU+ymPescsKYtZPH+V+iox
E8e7RB12DHQATwO1e9cQQqlGvf6VYWrpC3SssEaAvZIzYB2wH7YlxUxzyOaSsUY5
DciuYDQ1MuH/HLJZ3BT1NsZG5IY0t+QPYXFBEK3YtPQjD7BKwUaaXpBKO+H+K7VJ
jjCDJfQGSKo/zRsN+bzlSSEap6+Whj8Kihg9JdRVGMnb3PFqHd0Qgix11zvSDFRU
OQ0HGlVZSbpVvS6UbOH35XZUEvHYoTyaQ3qHnctdEa+qMD+smQk8LpsyZHjN8IrQ
QUXbdLsgVIla6QmyrwlTM3i/QKoSBRUKvP4Y4on/lzFaciBmK0O37/MnuJKoRjFX
HtBI2QiVHRkYJA6ltioCCcQJkvIsx2sXTxKeTIwAAF1l+oI2F7J5L6uaRAXX7el0
WzxZ3+3wYPt43MqrmaQVxplrlCo5vyExPm/2Z9drGjFUoc72SICUo2kQX/ArkpDW
fvC/kgfreNnBaW0LQTDUFTwgbv+cb1z2CvXBUs78dTZ7rbIp1/E4x/xo09ZvnWJm
G1kYLkexkN1posbd42cxkQ3+mk2fGFQv2kwmRDzx7xmBXuJXJ0kYoMBtWyPnMh1m
ztmXym4Z/HGnE/C95tZoVvkAbLUHlI9faf2+ViRXmQ7477JMdw6MPR/XNNeaT8Hn
1XgfiQba50R/p9eLjhT4Gge78vk2n/ryaIi39d8wvHu9129CUWGhbiR9M439MVgU
1E7zdBcTtILFX1J/k8xOkE3P40v1fm5EEgFrKIN50HknWjYYCuV4qcLB6akKjdvz
bqY5WU7vKT3rjYpKXPIfFDp2Kf2IDjSeQvxzTrChkQaTH6nu+j4S4bjyTKPK2MUB
t96rnhdtoiiEUtt7FSvCzjSXRu/jmvrG3F06V/URYY8w8MJiBwfZcJwrCL9KSsZy
41iA0V0I4YzCPLExOkxtl+1UcP/ixmt0tC4a/SgsR7F4fCBZgaf25ekRGdTAQHQm
85GqnNF3gdnTw1YMKcQNg8VQzB0Snd+qOltLhEIbqMNclnL4u+g9hoRm8qAUJXa4
yyyixfBCE4zgOns2SczOSWaE8ETIE/0rWZEs9p87+5DkZV/PDqeQjxwMgQ1spDJW
fwoimV7rGVpl5WiJKTMWaa5kOjnNr+Q0OOIj8jZdz0J+d3JCXoV2FKNKpWBLOcyZ
ev9gC4kPw6o2YNvojdfoe2L+w6ctz0dvOZYOX4x39U/1GSFdEq8r8WYV/qHjw9Xw
Hb8EceHquux7GrEFyGzrsaezLqqzvHpegdrZu9KVBLWWS7tkYZ6rR6yMy4yixLzj
HRw9/pZLkWPaJ9MWcO8PI/wuTbFh9Rvo931Tpj0hsk0zU8XuzuiBxW1GZdB4pJUQ
mFYCWv/pv5isytUWPkcUaG9J0R1/9/oostKRT8BhX6ZrDPcGQo5UDTJMwDFvB426
Xrbw1FAYaZHEN/urNNVGymP03iNo0t479mi9icZj7GAxeyzvVB2dvyU1QQtUJMUs
GbKMk3PeVsW4afl74nSoolYUcCIPkDt0V/YC3A1E8WgVUabRG0Cx7AW+rqYw6397
PaJIAsZKhkXIZP368dil7a8CebaGcCVY8ZlATRyacZQ6IKem4IJuJd5cWab48p1n
wCgOttJoNlDnUExakdDlETvWvFz//9Bj4jkFhRu5jQZpHB0OaX3dnR7twIYa2TyN
ftBqKA3LtayFfAfwRyTCVw+delwIVEf/IYc3fn1z4KdhHEae7yemDBJrcCJQnByv
sjka1WOBxPGh5KMLn9ydXaxREuX0mscEUfiMEGXe1YqnJosLV73u9slbu06mMSYi
Wn8lHtA1Re8M+7XeZQnDZ89WvSRp2fGkeLf3XADZn0j/ZWP9aux8elokgVpQDXvo
C+q+v5gYTzvR0WyfTypFeWnIANTUQM++PggY/dDjmGkOqeNlcBEcJ3d7CHPc898r
OhsqtjOZxjpVFVSWB7QYc6Svh3JkXob9qVzQH00se/81eGGBu0bsZvzVIgtt1jPb
/jhFv+hrq59jmOhUKGzfCW+R4h2z+K1NadN52sSFmb7K+IBKjYTR9vYOo9K6iZ4f
Qj4grra9LBEwyvLjBclTA7PXmUsXW8W0D46jVKR58DW1pI7CVpXaMM18VFfBZH3t
h+OVyiis8h0SQ1EkXfZU1Fc/IWgcg7EVeLYIKxgsue1QwtzytXHtNkRYXYXHKG7H
ivzaUvlQsRBjlmGL3DhM9MnYsVR85XJFUD4IrZquAOPjOz/ivUoFf2EFWzsYmf1x
sR5zS4bK0SyAOL3rmUZAS2jMs5IBfaPCfdeNbS1i8/Ku+ELW0TT1B6UYLy6FIlYw
mPP0OrHGAlyhF5OQeBHZn6aHrMh6Mk5cK2kJux1URCZEFMG73oYtgIUmhAK611NB
3lePSHdeKp3x5Bo/LD/0D9oDU1MqEe1W/+xm7J5KXCwKcXYL/2niQaDQPwThtZ9p
KlJ5DoXY2FWebwppnVBiFO+4NvWVeOc5j6rkoc4rQTnvdtpniOFjHdTf1mKnn2nL
Wi0w6XX7ze4dXZ6PAOVzS7gItkAYx+qW2xTA5ToHfHIsFhtVWYlGKZ5tYEij6bbx
jPTW8tbDxoUeAJjXLxhsA1stx6DtgIqp2uf4L+lqnfboKmAOOZcKWoHQ7z4xoi+z
XUuQNpEWQTTZ5j89Xun2r8AZOsAjE2JWRMXlxbGlPWljHuVcWZB5IwERGT6sisoh
ra413XT3wB0FIH6kQDm7oDB1wnlEWUvJ3mrMd+4oC7u2Qm077mSXT3mcqGoVzysf
SBks0F2Dz7tFXx8Z40FgecBhbQBp1XWKeBAYI2RW9+38dM4+Vr9dZYqPEuSNjz9H
CWsyRssagUtuNKrEsfTMdociemJ4IB4MBmgSAHcroi74812BDlT329k2OYZmjQd+
gV0/u/1kgcVbBt0yglYJuWn0DKXCcPGTyp/177ROxJMdVen61xX3AHWyKbIrpRXw
7SDNTAqyTW1wwinSqe+asanep9X8HXOUvwTYwzZ+G0//Ksbu3lhO8CjBfR1RaeDB
BDx/FCBZrB25AW7FqKDEF6f3wkO4WcIWEda1yqecpTO+NmfynBCEwE/+xzCbXlpe
vmi0lR5Q8C3Ccgj8vFlVQkLhq1xjg/oLzPs+QDoibDEDyyBg9CuA9cBPKg+9x2RT
Jjy6x0gR6tszV4n3x4T9aUjolH16ZAQxZlIGgZw1U0+bXH1QLI456A7dhtmGJnex
eH9LE97IOp0AmfeaKUzultM0hl5PjBr4+vW8ASxqn1WJ8EgvJ1SzZFIJnYiipLMI
VrXvSUSqUGkcDPd15x/28K83WzmQOaB0IKHwaTeGyfBa99Q+/2VIlft8k/LLpAYJ
SbxAUa+eFEEwJv08YjPGClxi82mjCmitZamzhIAM/mH1TPdfxsmpZP1sroQr39hn
BM9YEVSIRUQMenkww02tx2Mt1TtycjT6+3qKDkSWtYf36pJxBuQWtzIj4HgnoFAj
ZBAvx6GzEEvdACucgI29ITKAHaUFlrRbvN1u00r+AS3u6Dcfn4jED44pqLlD82F2
tyFn6BInLmNZHSguctArHlIupcqdVIDtH5JZHHX99RNNQwFkfsEjL0LiqGnM5+vE
aoJr0E9Wk3bL93D6XkpelB5WwPecdbSMWhrUPuuiAatZUDFUtCFZpN7H4SGhk97w
cyLAgIcffEw6igXKp3fwgUOHDpku7TrZzDiz8kM/BtQaZUnnH+6xaGVlHW1hwSiy
cw4S1PGg0YemcoLoxgOCXeRCPFNFEFlYU566V+6ypAUKu3YfwAhnRFhV4PqvaXqL
T7xxIO5VyWTvolpA8lVOyAfxZZt03emgQ9Mnnkr8EGsOMBS6ViHjJYoJx/K7yLjA
Rvil03ap+7aVs9TCGSeza22ZPj1O5Li76R+bmwCb+v1BwPhWVoCU5p1wjkIvklnv
fXGbKb9v8tYnA0IRHSCc+LgBPNiBbKobGaAjOmFieoTvWV2Pi5CuX0BFpn2bFKC/
FS8iUbnuP2QCxFdvBTG1mLINfDFzlzXXfkAQCtY8hwRuSa7QYu+l/usOQd29pGR/
fNN2RBPmEEVZODtsRboy2Oj8KnRVPSgAuZvZUb9Rl5THYf8kwK2xBsvQ+BPm4W14
ibTf2oTA24Nw8AvYFrG+iIQ2JchJ18SWl9neGO8SqhmsDYlQQBlfaLQ10oTfunxj
iEO6hX9Z+bedGAwbLYQr0uz6ub7afDkiyhIycKGrCN3FKdeZqRppM0pFKhb/HjYh
ZhzaG9pgFBIrywKqgeLP3rNs9ZzzCc6Brr4wFiQ6JRbRE9pLcCLt3/xU2HBdPtYF
S/ODWC5HtLFFZHByk5BCPVYvtFxrki55rImKHayEZ5tlL60QZoqOqFlPpQ5nwLA3
zcqY+e7OGOJ8Wh9DybsPRhNuDkgav6HPCB+Qo99QPnl2NUVTZz/GAygruHU7NV3m
3d1qLHFAKi+5//j3+8YV2RM3N99wfDcBrphFqiYOarY/6iQR7fUkFXK18jN3w81f
2XQh6+ZKSkvWEW5rmx9eVJiLe1Z2DupmoiqWpTtVxWApb/Jk7A+HJWZfULm7cc60
kbz3SnJC3KrUIvyUHbLIQcPw4K3hlgl47yZSKiQyXxWPM38Q2xaLfiKzzXqNNW25
ody7hW7uxxpBvsFk+kYBV0tpdWND6lf9ny4EibZ3vcjptSLQDNYXnVqXEG+ZnZnF
uLxR5NzQXCGFWDAlS/70CbIUmO3bJuhsAnS040vlKpOAq+hc4l+eEvuPlqzqmtZ2
ha+5vDaqyy1j8bw+Q4M2j6sRrExXFQ8EjBPT3eRqr0p3F48ZnhZPFbitDCdMgtCv
CVOuGI13kUrXrOqD/ZShXoCnNnzFDgTpgyUj/YP0JH7jnMVFd8/fdow9C1ZZSt1i
LRtffiN7mfaOvKvVfvfaNlcT0sVBR6WS65LpAtNWoYMOh8Ez0f5CDeJ4I1BNdT6+
xw9M7GfJ1zJKRz5TQLt+dT832qVRUUU2SgkI6/PHLLpQzJCCoXeGZ/BOgGvFRh1/
1zZEOwvG2HhHEYE2AfmzBehd/nv009hlf0E19I/pj2Stf8CaTWdUGbCMbZr85mm7
QslAAytbRAi4Ko8jpbB0g73WDhnr9jrYzm/EkQiczZ5uYHs10v64CT3AZRbSZ4nd
PRUlZUxGdkJku/2JkoQ/PrHNG9ptEJhkGWZr4eruRbYMulAqjleO5lr8my6arXrO
qtvia05IOT+x+CkDcc9ZI0dzMBvTxpr+o0ue7ykfjRuZgxQDlfwn7ZpFeL1omRZS
bH8NNV0idFTXdhnokYcywpTvz+cr6WrW6bq84hWOLMOsBObtQXRf7KkNVIDQYrI6
Zcvuet+yQUFHQ+QBrhfxfT16tLpGHI8amdWqt3IAMJViuwmXii1CJhtz7iGf3gNZ
jl4N7SswYxOq3e5NS4c7xto/nrK/3tIT5VrfHNBABurq88Qc9UdV4MeZyePIz2Mz
9aVrZFH5sTWKRjUOs5RoUw/cAys0n/YJ0klhSAQekpXMt9EtMdq7150BF96w4V9N
TRig5/lZ8HoCvEGFD77TAwg4DCkAYylDU++bJjQv2mYDEE8FNbzu/CY8VroQD/NW
4xR6gfZM8ahp5wnAVl2fEYmvicBiOUyUbQMHL+ZIxrUcOd109iRX0c51JBgGIO5u
/J3LDd0wcedquIUjLrh3EvVPFCx4mheFRtDwGvxURHA1I7cvjRAFgaYvK8KP2+o5
Z91tVjQ3uY9XYa9r9oqpJmZx3ftj+bBA69vPjBUwcjmIQ8zLi68iR4VIAVMT751g
QkOEddxpUU30F+k6Iupqu67Je8zBMQKJR6KcqKN1JJwFxSqz0hwHD1mDrjLTYx9s
fhzTNP5YKkur1Gbhi2S4QmdNd/zrEeUzpPbdxEYWnP1ZFQOnPM+1Q+pjZs6fTppG
/uZ8SoSDruk4UXTaizCLWeFKvXX9byLkS9ZZMdp+AQ/4ua803rjk6iEUqqO0fTMy
821AJCZnZuWr4UtVQ2C8wspFvfZRmxSZz2R3Rmj7CJmvnYXvbDaCwXWe961kMOhG
t9RlTPEptOecewemECdY61sb/+azSJTbzOCAAulZ2Q8W5AYoF6RdW/qOwU1QMxQa
W6TLP+5YxthfXo/NPWQfusb/s1tpD5bCgrxfkn3LihxnyJlYsXlPRpbDhZ/9D8DW
k3tegmZuNhDoMyu2jneA78xcJcgaF3SfmtKhJs86LMUGmPyn9rqxbiXsgiGiw/Vy
u8fGd86vDEFgD5MdvoOzx9+CiKfuTOk3rBSsxAny/MDh4O28CheFBpXYah7duM+p
0dUSy6rUp/qctEyCjTRNZSOQA8v0H5U5z9BjsG+YWHcJEJv32rW0hS5ux5T9wq+6
vW5GTn2+AUW9uH60Uz6EJD1GeA8yKfKClPg6Yyoe9nHKUNIzus1T/zlQoN2V1wtH
ZFefIsaK8VMh1Bta0YrCXsSeIW9djmpdiRle8DDxIiDqbyGn3a1ECDk5vuKiqz7K
yn29UsJjTyHjnOdfkD0Yy2Ph6xpSt+vzUvR+dQAZPfdJi56yGriEHDFdZCPGh4kJ
Y1M9JnUy+mkoWKv5n7EZCoSF+K1bVm9y/6jxI+YOz4EY0YGCRUWD95EVGE4lGm74
HxmlJVslnQi/5qsswXe6X8TyM8XkI2Mbd0Ba4cxwnLQhQXqL3Lr0O15x8BnPbbOW
DsisYAvHV7XPaDK9Ae/DflIwCbeXCfzd2nZ5+o+0oe5jDvIvugRq3JgpUVo6k7Ml
qrQrpAwq1JNv3HmOyqE/mm/COShQ3DajqKRpzWQzeuEe+uJ0YL5GaI6WAM9cvuhq
3d3uXZu5yLYXCySXcE4lu2XVr3x496CO/uTNG1wb/u3LGiFgZlMaQelNGMM2NU6Q
vAxst1g82gSjW+C6al5/EYx/9pqlOPiQQ9910NP2b9gteFXSa1Aa51pp1VZLmgha
JEg/7cqss2xOeN05WaCeU1Sf6jCtfFIAqqHnGBc+Ab/fVTFwXYmi+rpOPtl0f8VZ
4+pj53NMsXmpCvxupBkw7xgVqaYhhVNjY1zd/KQhbZ/RRNBOHRgbA0NiCwjYW4Mc
NomFm6msiJHK4wgrzByySH2XDdGrRM4ACXkXc28X2ydEFmHSPMQ9+sGsj5bgRZ/w
5iBmWHRus0XSP16m6CeCSrtlQ63LFZPpymX0hr9X12nc1jJ1yEIrD27QbPdjlxeN
nhMvL9F9tLdaLo80y845MWCJJU1CHhLBlp/ZIuVv0vBT3LyklLvjIe9uc2y3qAM5
gGgl7rjgnDNChZ3wCqClcTfn4spT0FUuqcE05WSnC7D6u9JErUGMdsWR53KeukPp
UH1Lk2ljDaIuQZCutEb6Q2s9bxw3EG7ucyCho0eHSYTgHwALbQhzMOkeddRRys+D
63H2aFM2oU3K6fXxsjm0EDfmo7nzkaE8zM3IEwPm7EwxNduPNNNGz5UCm+H9qTFe
jpCubEMaseR6iQMOdxsx+G4k4U2yJQ5k52xCLaVhjYu4m0Q0IV/1OqiOm4dMXBa+
PZWVn2ASpTwH8oL534gjey/GuTn6t9NHlyNbw07RAagVbOVbmO2FBA3YZw/08v9I
UfO60c/pXQiYF0ar8+IVQjfWdhyek2qySV4QM7v3cwdHYYkbrwFJH5dS8DpxrxFn
0x85tkuBGBUe6hzdzcgyhzYc2JL9Mc8caXHWbE1uB3lQp8l+WXUHlH2h/Y0+eVzt
QK/J1WWec5tJ6bsCBdo8mCtW60qbeGDVzTNGAwbN8GMP2819psvKr2ih4vewju3k
BGakB5mgcfSDa6OxO3Ooe2d1bF5ybFoinAB/rj33cVxzD7yhC5EXnTu6BosFgpQl
oa7yyBrBj/q2LT+70fk5nHN7U5IY0IXCdFs40hDbCEiGYOSCEkfzAseyZsn7D/TY
pG/zp0Ff8m9sDBEGK54yC7GhOl8Y4ApRCYMgCRnce4lQPIRUfXzCrtK1VJEPHVch
uSrsJf9Hq/VKIsJNIN9ujxuHba4I9yyVSsJYaECSlyPfgeX8OL03vxyMGUbgsKOm
1gj1/X53mJFaZVlxXJ/S4NOdP6S6Oa8+HBDriAyY2VDN7azmZdAIwBZTiSX4Six0
p4LnEy9FyEmsKUVwak7Jc7PKqvtNJbjjbpTVapGzVCQIioXuv3oP+oyRkskNG1rd
I+kUHQ1YfzY6GXmXjWU5PNY6WwVIZPPrAE+8c2tCil0V+ppWIEZ96kvbjt7y/7M6
0KqIDI1GEVa4PGnv7CjBqCQzlmJ6A63my07dKx23BO/WgilPnpw2lZtSmR+90s4j
xrHwo/7ssmSdefZv1aegsKV0dCSfxWaTT9yVsYNlmejo2xlNkrLp6utmGLtaeJPs
kQ8la0nUWyTYAqZII+na8Ry7zPqP84cIdX5T/R4eDmyetT49OkAo5Smq5KH+bakp
NbJXEPMPxtVAAgavwhM1zmSpO2bg34tunIDBLYUr8nwdRpugm4otVqEJbqbrK8WT
TENhqvvMhvjLnJOEQPb1DRg/CD2uW9I1FXJLicHbmUVD/qMH2k8CejGIUp7uhgR+
Sm/yJLlaqnD9jOgahM0qR57vQvBWLqQMWLp7Fjy4HA3/j2D3791N5yok/5hHh3kY
pmXrjWXvofkxsC2I9jA+GePKVjLUYYsp6HicA9eWWs/o4d+CeDuB1kLs6dzVRQSc
gIpSwr1fZV6mK0qtQLaN8tpMnxbCPbxTRPfrJysydqcqg50tJR7pgw/7PhVLtCLG
ZuPLFlwCuEzLZ9IuplxJh+5ExDeR1fK47HIQUNs8sRFOrfNWz57mUtLyl65bbElm
x0tGp87qAxhwbtWKA5MFCmc3dHLxK6N8MUArjn12AirC83AKAg3avq32PH2QPwns
6HQi5M3+ulBz0XpLDxJG4MO2WV1UYvrPxsMQVZOtkUr2qyH67DFrChzdx6d1ru4k
DYnVr8I9EFf8ITss7gESKwsJt9tMGXZ2/2RTtwPfOW4NE+x4BlFDMlZlArRrtemQ
FpE591G7laVZX4xJGYJYTAr7ZWVSKGxo0GZ595JXxe2DDzGHJzPAAl0vaWq05Wvl
Y8kP9xxU+VbXypNMtXmhGyC0ehxXB+MnoZeHjcilcjWbLRLN3wrf6kj9xNy+wVC5
09zot+8gNSNELBfUrm07n7MBtLjDMRA8xMS9rNKKJ4NGrZ+L+YRk+4wTQ4SPz2UO
b2lcEo/VhHMdygvMIcJhs9xFZtOOI6fhFE6RPLEKxiMGNYzKbPw6Ox/xLc8LlHk8
UQiRBI28FxSdkGIMjzuzbzFlt0kZ/rBwLoD7Yh2ZNPqg8blHvqYeWiKQbha6RYSG
hZSP/AT6W6cgCDAR1oXdTId5VAL8bM2wdgU0mKpvh/O6tuxkCF/VjVvJhRWeKaB8
szRBBOxlEN/W+5RNOF7oT7eth0sSn5D4ls8MjNhxksf3MAlyQyAunaozqEpVagqu
+XselmqbbxfAWnCRBokQ5r2K0O5h3sUySefp1kgU1qT8RntVF9nW/x5oSVK5e8Ty
KoCWQdhvte5Ccskcyt7g0+royCcmWkisAWtrH6elRNxAijKemR7oKQpTGtPEdMdB
SNc5Z6LlmTXCMC7301jz1cXCMN5OWqhqi4PmVNXY5zPHr+1kCpNXKJKkUz3mk2xz
Hq52aRn7JMrwUXEisar+5WI3aJHl5kGx9JHC3PCVeG77ZVVCK3pj4U1hPThQHL9g
YorHucRIVprzu37Tu7BiEfYqbfgtMEXTuNtvRvILhLA0lOlZzQlguz7NSylKrWX+
yklLvA5WTuPEIUzh/cEEtTQbuzhmoJgAtL1ETYVBI4pYerdkQ8g8psYwvYjpWQ8D
M1zE5QO/SVDPLJBR+mrQy0VaqzjJDKAApaNRi/6CToQ5eGAFByZEwhx0WK3KnVGZ
T0laLxKvptH92HcPPXYYfyuyFXrLopc9VJu92Eu6ZKVK/mqnqpZWe+H9u6WMHm/v
GCO7G1luQcdoj+kmjhfRBsXESqDSAnyftSFjeWHf7hjUa+eJTFk4/t73yGZ9Ey0/
Z2w8cUXwwxFWuQZejRqwfBd+h1wc5bemS187Nzl4ox/fWU0jRePugnjyQ3MP15zi
AksUjp7S9Dy9r7/myPK//goaNxINPsLxWSb0VuWzr2ijdZrrkdZFCi3zoiJX1t+W
SKqCLNwjl0/wJmaAJ+hMS73mFaDpeSl9XyaPckjMtZ+eVyAtTr28yDzbggWhjK0O
xQtpND3vDUGW/o52yQtrQQD41cV2bekW8Ac47v9zAsZsGb/espBlizqwNoskp5+v
8495U+o3Rh3Ft63HOR+MM5Wt+ndC3beL52TgWr7TcfSqvWZgxs6ZFCggQocuoUaz
lOs/sNsnFnLA9/rm+y1fME3U05Fg/kWB3zf6Utx/n2FfN3Nxy6bCTHepxlS/qSx+
S3S/RK/7Fy+j6P1aKpBDq2KIqNCyg2ODYZRqR5gLBRBN3ADx5QhKemTzppDQSLFI
nGy7s8qSgc19UlaW0Txvg/3s79z553qbbPTHChnQGy877tZzFKoSsVFgpFN4lUcT
2lk2ssuHB/oxbcTZWfN6PrcAcCbB6XHonO+YOpZT5ghOI0bYVEtO1S4TgupGaHfa
IlbxlTSKqxkgybp6jl5udmwHpZp25zr08DAiKe0UmlbURahZv6PpwgDy8+B75iI5
IJhG7tHtTwPCfuPs05c4H+PJjGX+fSGhUp8URNAkVCHEkv6VkHaqsQa+ycT1Hx40
kMtuZIA/Ouj2TQUiQISUf66SnAkE/reQosBNUDeIHto2f/0UpQfJkRXzB+1Hqbep
fuv7usrjqAg+c6M24LrjHyWt5x0k8ER51rjcFdZUQpFEinmptrt6W12AxiKsRsYu
YPjlJFUi6UqlAGutrYxNmxMsQYNpaBeD/YtkbAN88LIUZoz2gtnwNhVcPL6N6ivZ
dowrnii5tfJtN8IqCNXQdInlBLnmJezQ+eel0aBFq5zHEm2+1TGcIe9DaFk9tm/z
rfC3+yuAFoOEEHX2oywGFsqJtgwoMMHuOuOjvLesJNLKOrJIKYWybejjDL4OxdSm
aWe5eKqncwuvOE1LRIPkplzpcp1zGbrY+vJSCebd0YNIytMYtUO6Qe5QA75hREUE
wXYdpNZnifQMXn/00TyoecwByMP103v4GLxMqu5+aw44Qofj6PMgVBCjncGsWJQa
hFKrftLwmfRV8vzo7UHXROHgrayCriI5nniGU14uul1vBOfKLuUEidKfnk87l9Fi
SWoOYmsnqJGJFXSboInFN+voUOo68qXz7syrdisEnYleJM396fDdKOsckvgFJsYW
9ewkRVQLiFWa2oxRWtf2H1sXJrqTqK90KGGprjWK5djm6Gd0E/QkiFdGIduJ5NnR
9V/chlma+H//CnhMjLh5H+AKR5aFIxBJkvPEp66Li1jSgDvp4mnQ7JayYicrMpD9
fr9s3ASkRTQ82T4StrDIv1u6P2N+f1zlUT4CWAokStXTWQm2z0CZ3Nx34jDKjCbI
gyk13aUh1kFA2A6J3MjWe9SEMaOC+SG3YZP12dZjJzrcESdtTRrQ0no76EDkM4x0
4V3YUBfAxWbklzWSQa1TZ/foREaVuJVCPTgNsyWafknjYfbKkqD3pL/XjtJ9BWUS
sM4a4mvVyc2Ri+SYCuKGaHu/GafO8mlzuIWl86RQjBm/ZZC1fDLlQ784ZrZFKSBj
Jtfk/X7KMi/V7eXndd3XyEOUhMhXpZyWymw/5H69Qkasm92DmJbHuycM9oURcn8c
Pzlz7x13Yy1UfFQnK4asGkboc1zrLLWGfw/eAMn4bmN0ZIfynJP8CyRlkjk1Gqxz
qc+TkABFEcxLSwuo/KqPPjt7hQ7irUrXyUU5biu2UNgJwD+rBGt9SEn+pBduiXyv
xzZLHYy4V1GDIpTQEr26iyp/P4oeWkhDuVUhREHZ6VnV6vWcgdetbyWGYEhTVAuS
sGlczteCjJABZvwpISqMUBMcs6muc0f9Hd6HdIGmTouCfX4z3BrQO90F8+Fz0i9g
YV4iyRoPWGI2E8z3AavsbT7iRbjSVD7e1jtDSdOK5NkmJ4f5cK5lmXI1f7v3iAqr
cSIEx9C89nflo1wTM2YfjgTEwIodvUdy1N6ThqIV6eQLeo5VxAR0IEBL7+GPSCXP
HNSsUw08Oq39s2jTbFlv1ZksMpBcWYc/aJKJN2x2MDzoOCriqqP6aFB9VC8mbe+x
0YikRuYqfiDscHZ+de9S1xt13i3GTA5T9v0mLOERtXyb/QV0DN3MbRSLLx3nBEeG
1R0dxrINfYznkA/SOAWhJS+gUDFwCD53dO9zEIWIQQLjuEy5ZKklZal65O9ygxQZ
9tOSVPxikbLaBZBpjiYUvyneTZl5CUpH/nxlBd2EXqnD8C69VA7gSVsEQtAgl8K8
ZLIQtHuRjXFu+drqMUO7K5VdUemFcpiMTpL45s7L3DA+Dqo42SoyjMsDJ7n8sQAj
0viDX4XmWfbIpQMeIP3FfvviWVJnmaInzcfdlt1elUWKA35dir2+i6QYviNOaVKT
0fsDT+sy1OITaTm885gvq13vodIpu9ah6LtUMAovYlMqrrdFeVmm1cKURmp7UMQe
CicBV9VUXgJZkumxVnipbaROnFYBNWFv83JuGONeQq4439YiG/zNLjOqzv0hXaBX
VAwy4gdzydCUQ3NPLLuJglpc0b8c2JHbH8p1rFyM2Fkc3IPlEYc1keqHFvmXsZ9P
GwwhBcd/TUxvUJTMGrlQa28wH46BAFloFGK1TPhQVoCK+S2phL0AkadOY7SirneM
hyshEn77vfEJI5lvyGh1IQEBorClhe+ahFviGs+FdoeYLy4KIoGFsoGoMwiRi/sq
gzsBhbjySpujE4kFn/3u4ZceCB7Zr518He5fNK1KLE7X6zv0vUMv7RHHOBb8iuVM
YsLmbZUDanCHUo6JnlWAiIuQrzPgSqnF+hARZ8j8gHuyATOAbVA49uIaj/55QfTY
QkGxhf8PEqnSmB/3ot/VhmR/ljVRhqGvi9s1C5kROM+oI656x+vJNTj/rHkkRjjS
lFHiIdTcNPNGfm7C7E8ghDcrkIWus/durc+nbVC0fgerZFYLwLjGpU84p+gCf7+g
IWcI4qxcC+roPRek0uDpXd9QpjUuXcZR8aOwpUh/9TQfYg4YmBKs9yg1UhX8Im9+
9zqephD5StXmYz7fPcqkD5Fuh96ztnqkBCmCTiOda+dp+90Ec/QvOgZKufmhA4Wc
0h5v24RqgANPa8bn/QszotgNCJOyocvVJrV7S1CQ4+6ZQlOax8wxwQDn8EYdMNNj
Vw8rd4r4vr+j2ZTMK7cdmWRYpXG5U2sXGxBTJSdme8njZwQZv1KPOVk4Q93Y4pkM
iw8ZwWDT/7cISI2YZlcXuewGYDl6nFJDd+YbldEtS9VCG2Gq2aVUZA7y5Np6EH0D
A3hMKAVaeBo0sQ3WJfOQQEmUItjyqFzmcOxDvOOkyGMFlwTrou/bGd9LQTjbKPgf
fVs+pazqewH+uWidw6KAFh9VnWTmEKqshFzjHqGGphKe875zKrZcY+rPwFjoKxrm
Ht5EfN5ZUH7FYzPexATWtinNyijLTw2hvLxDCLqkkeQH3ncPS5X1yWcbEx1u8ivs
hn+5I+jkKEbbhGo7GD6llgOuGWL5tWZ2A4Ql9Or70nPJw+N5wSdoRvl5lVRWOlOA
9LiEKlAlbAeBzVptT1gVGCTEX9npH4xEVb9VI4R0SPSu7EiI4yXYUqBQXnd9TNGD
u18OJjTzh9VKJQihqOf/NyT2eeVA1jhrJ4Ldjo3Qkz9mDup5m6darKG7Zb68RlDb
2qdXkLMk0Ankz4sej35Zt/D+W8vuanF/90iod2MMtjZkbmRX6qRFxu7MSW3G19rn
PlDUbDCa1U3tb8GQzqbnj4EPhqXIWMfoX9a5EirJYI94XhS+p4IjZeFUTaSWH7nV
+D2OL4yP0yvFilgJ/EdfIeHWAH4RxswYiIbceE6+sWv5jUGoIF06TC6rIDvqWGC4
OQkPDWI+xoQ6e3swjOTjEZA0jZC3MnClhIQRs5nMvasgUkK+i7mZ+xr+nEU/pLVV
6mqJMnlzno13c1mJnUwcesqg/xOIHBVs0gxPaOP3/I2j4FuRKzFI6G8qO8wM6Pus
w0ILQOGj+M06LCsm3M63zeamBJCEkNlbfcbsGcNInYw/ZiHNe7m8XLhflafCJhAJ
ebgr2f+vYpxnUWDMwskGeMbtt1nId/RbSyrvZrx48MrP9srWHssosN572+qHr9Hy
mBw0NacGHDKPw3QqUODeWdAZJo+7G9BB/TZ/YOpWY3hfLPTX5PahcGU0UNItnitQ
U9R6zJxXedvCzq/+9IA62Mt2Fouf4uXUFjPvbnWTIxm+iCFZWpfMAldT4ReHisJm
90R2rW3gB/RGxnmVRqOTNQBO2S36y8T/G0+GLEtRVpGv+GguZmhYXa6vP6HwGKGr
MNVo5BSSxxj2qqyJRKF8ww6F51QoJ1FoMB3Kkdszl6cKXuubK6KZUT5EhRyhNzn8
tIKU6XFYYExNKB/4vXhslk3PYs+ohCWyQRFTrCgj0OLXa/GfYfi0DiA7kvK40kQz
i/+FQIG56jC6fjRcNyIuTIjHrQICCksGvTgLzh0ObTAk9bWGoqfxOw0j4uyEa+FE
2B+xlZHZd3IClEfBBt0v0bgrDsRkcDtr3F8KalY03ukqh25FL2qkBKVi3Y8qr+00
lw9f4ZkeJMZmCprF9SipztAQ8sZh9mYuz/VkDTNc+lZfRW6Fk54xZ7zVK41nJY48
wv72H/7eazJM/P2u0UXtu6w3V2KN1w/71gfUpDerp3BKMrBgFa1Ifb4lBGm6b41b
SdLKpJmZpPdPRnxCvHYo/ManxoZKcXegJAmKQ5Ywo8WSt8WME0cacC0AyDZnI6tG
YwoLKCy0CxrI5QDL80ugL59Bhh3zatKQfWhYNFl6QhS+QUjdlaojWDO8R0GjiSFA
BlDBDkhJZ1l+JOPSINoORgEksF9LPQ+/qSJbthG9ZpJwXzVsoBfp+ZeXIhpNfyi8
pcZSHxCL5CEeFqSdLXhsALEUsDsaFuprJUTnmseZZqx0GmCbUgc+UWBdfyrrm3ul
wBTNndXruFFidJiSbuX6GX1U1ZdIMxIfK61b+WqIVFNHHi3TkwNB4kWZDfDgs4EC
1hY6VCNQ0lBehoTQAVApZp1vCWVO190pZhDyZG1N3zpYA6XxnNu/N9f6DKkN07al
O7wcIFfzw9aCWNEsrdsuXg3XFvgDSXZ1dGlB586GPbx/dVs0bgmlBXh/79xCvFf7
0/FDazjERaNX3k3Yanifu4iUbylfLFI39Q6Oi78SxrdsHaFP5klvUOl8ZIPncDEH
hLYNqymFe2HU3x5xQTaur/gDN87WU2uBETf4tzdrHRdqZe6q+Bf+PSq7bVWbra2v
ErscaXuTpChpbpZ4fnzLoYu61/Rs2DkHk/Iz09agCB5pvvidV6KePq9fHt1LQoDY
zYDKbf3u50/7nbnJOu9F6p/PuhAH1xcstizpSNhT6D1Rc+nvEzQoYqcIi/1e/d9L
4No3/UC249+kD7ndSGiASqr4CXndrz2y/lLI9lbOOX09FjtqnCoWMVLXu4xsG7ZC
L/J+9NXMDLnYR4e3ElDGF1KpQcT9ICU7PgVMS2Uimber8lyNvANm8cn3g9OCUHpe
hwDjsA8WaXhzM+THbOfOru+OuWagdsJfY/eB272ybo+8ix1SF4gZpZ0Q1tcWkFl7
NnvJPGolIIAeY3akQv7jhPqkdb+xieIC0Qx2wnaETX02roydhLcLiijNI+TW++qG
eUhLZdg3kIAsLej5l09QUX8GfaxuSstlXxVgsXlUmuhkA7xJi/TGi831jIgWbITf
xy2/lq07rGjgLcSGolSaq87cvbiw2aEeeitDVqxZeYYh+JjLDMYCR9UpX/qJCo5h
8UnsE1tT3Smn/XL1gguYAC1bbAA1FvfTfNeA8bRsINQnwYZafPsf6KRBoV54+xy+
0jlfEk2dz4bIXxJSWNXSoHZtzG9UnsPbzkV8oTqxEsqGbuF52jQNyqTlEkw0T1J9
A3+UqTOQlHvyRU7+ZvDkNjgfQ5Y/1MJD3okGjKi1/KFVJbmXsNPhD3Ll6c/uk1iq
NP/2Q83iHFwHoDaSVsGsBN520Ab9kfzD+dxmKgXKYOePuKPNGnZOnEUstgZbKo75
LwMJezleyuPb21g35tlh3yjap9XIpv3sPuGkjgxdKNqIEOOlRaSRQ9eSe+T2e1B/
eVhePHM9QrWRiyHBhkvPX6NfV0R/K32GRNI2+joMW/CgBLaA5tHSDJ4757W4qq1t
a2DbUcsU51EjHc0gvJtWfNkZsWfd6HZw8VLtXqk61Ejfa5MeLU74DUauxNt+CS8y
WfR4khNA/iug5pCB+8yBO1YiRV0HeVV1sXwVKemdSGMSmQ0v4+mljE5ZcugdvbBF
lwFQyJLFbg/oPE4YtlumvPY7lUbJFaEuCtVIRMeujuZ/cZF+V5rmgniZpRFh7hx+
nVqeGG36kNhKfymCRF5rgdTIxWD21EQSUmymTTv4d5a0YQoGQJXxGnJe+zj1A0uv
wRUbQ/fdnS3f3G0PqedyJ+jgfNka9AdbUO92vgqeFC0D1xq/afw8cL9Y7ISSLJhI
FNo4ocnMNmHLd7XuchDtwuMFhiN2hZ+231Kmta0QjshCrqY8fsrudp657WPKnJ+h
UxF+B7P/urAdfjS5SgmKPRLjOdmxkJhksXENaQ+kEFEwdTpiESDeP0ZaB8Ttw+XY
G41tpNIWrVjeVc1aStni2XcH/UX9JL0yrDdVQxKmKsCDZhz7/dAAqJysKpxfuTej
CuJdn9Pjnl1FiCeqZLlEnW6WowyOZ53z+4jSEiHmRsJH612qj+NEfxaWaji+Hd7m
vmPbs84FOTbOCtX4LEKGPbRRyDmJ6ulDUTgBmTpu9jXngxTEm2AhYCpiXmAVgoE/
x9H1w/P5X9vo5/7owAockbj44C4DBSGmnK4h0Db4sggduy2d+oDFPN834M1y6vV8
EIGKIA7A/cKcmQLBH/P2z7gb+uoSXHatTgWhfCKOeadrAS7OKBl1psmtf0HWn1VN
H9s4cPcA+eu+VlfgANLHBlgQrijFMh/8Aa5M2c0VYDR6fCOhP+JgiSvozgKE+6Hx
Zt8XoKtEwLsr510i+mrqw2iU1xPj1FSTnOcxbRnzvoZ4+zmiwejXB8xSZfts6R9t
gw86n+huf4Osemkdf0toRKpZa4oQFywn2/lhMyqfhodgtqIzdsrhXs+aBOpv9orI
OTAdZ7LvTbZMUJAc7W2Naw8HlsApe+mokmBKtFw5Qt+OXzt73+tcQyA2ZFUWlNuf
AekxBoa8uRKFumvMj973Dovm+kVRHQ6WAvZdZxEpBxdZQmmwaZlEaJ6bA34ftJ9m
tXOmwvNCpQSzJkfR2Esr3S+i0Ib4/NZPd5cQxkcZxTuK1+eCy+Bj7fkXEmpteWzt
EDunyIr7EGbHuswnjsUN5B20gGsINy2EcmN29ayIxX0kDYa90k6wFPjyOqvrzF4C
29BinYnrkhLWcHQENuI7RthuLFk5qXo8zZCL77u2q0Gwpeg/AimrZinuJvobhZ8U
le9ZQ34LRImBtk1w7zNU9QNTmRw6zRMeWIgHjyEvfvE10uf4HPg/PwM3r5WkfIOa
l3Nl29mlVpWQcI0zmV9UTJypFWhbg1/NPJh/UK78hmXkNikOJRv4JKgkbfh7wdBo
/EFZ9QwM/oTRDxdQQ+mHIkm6oumsxZgxa3WF2RNmoFx2FLIWixD7mDg6P6b8oOz8
A0AsyTzZkpBUkJMAnVxGnbBfNod09oUOgjKiFmQGNPAYU1dLe79F0lzMq+otEZq2
RCpNGnW4g0w4oUXBPVYLTd0hMagwL8AIN0UI0tsUg4Hxrf4eapfLdyFlicmZc3na
VMS3uGfuglm5fDDJBJAuqBkz/Zl0iTW3/KbE/jvxpZgYIGRKWg0p+gQEbSb5U0jb
9zZ3i7sPx0oxh27X1EED3MpFI/2d/7VSQzyW1BHktkt6Ww+vG1RqNxnKxXh4hdWw
lBf4KfctwDd0CA+Bz6MSncRkADC5y1q2MFD3Bk17/ekd8cK/oknVO6eoGXq5DHPr
DV/IBlHraPgdGYQNeexU0rJ/259AovRGU2tX/o7Jw57c9MjR+4utmnbNSHUp3FPh
e0O9dLD0v5n5E9paU2mTjMJqDalhfabOyexmsSmBk88sY/IF0MBVeoo4zE7dDCHn
5rTCdDN5ntg2SM3ZTSLcQwRM7jZCNcQ0QC2Hg/XcnnPNIgnSZyCQ0khk1OcCU6Ni
JBVssFRFXDB+qBbZeoSzsPwCWGFlcG/JujkcxwpfWL15GYAnqWQaTXotKK1sp6qU
/8hj/kDYChvRzsoN/zdnAIyXYbJst7uyVQTk4kBHCqz8Xj3lk0YL/GX5um80cw5q
CySqXMQ6zW0Qav+HlyylhCK7iAC3aoYOciokZYHIayizJ5eDXANIsbrVG70Pk2UI
5Ml0Zv0BuY/jRgnp5vpX1j2PvnqnN8HoFlJ38+sGfEMXDH2EfClxH1eVwtvMvjnM
YNuPjDRamsjTOCdHvwF0poa0qATJGP9xtXUCUSH/C+hNfQq/mzJWP6fsN0RVEEAf
K1Oi2hWmEuQIne3uHbnV+166EqA/Fg2BUyT4MEjRy8wX2FwC5hXDKiU/6oPi3Ywf
N+W7UhSb/nK/0AKOL/rcvUT8zE0Ra0wsc5VERufZkA1Cp+Jb/5vG+M2HWqbB9SsL
pOLOBSAAVavx69kolCcb24Q/Ubg1ShupyHCUoShj8D+LzD7PoYlYTL4niX+ApUGu
5i7mJyssSl+8/5VEl8a4137BMdqNvy5K6GVeHFqVW2QO91o2U9z/ZEjABKBQ3vTZ
YBQ8vcV0SioDbr4GyO23xpRXXj2Is/GJddCb3YSqTkkaGwyDa6Z1RyEtGWRNDt6y
er3hCalGs+Gxnis+YjQsPiK+jfz8/y69FKDxX++irVGIuU3JoWYIwWngJIeq1ZsD
EuTKEW4RcBxHz7Vl/QVZIh0JlZ6Xg+JGVKDAsdBZRRC697wQKhDTviAPFc6YUrEL
sEldPlHsekU/0BvVOhjcHTfYF/3SWCO8YSTW5Nw3BewK7feeshIlI6YqHj2wvqvl
lyS07FGDNkqaJBN78gH0s3dgpFVif6Q2nrvlBx23tB62r/US2d5YPpkqcEXmxo/4
QuG6Pn5LWVy/pUOLVngUISr4XM3Xr8JjthUDcEb5FDVgeGlaPrRP5GgFgwNWhaUD
+wOfUS2mRzJgf7wVHpAQxCry0QRiZjLvhLuZnov8EOw57rs35U5jyK4i8pcqW0L9
odgIID/XhBErhmYrHIoe5ZtJP4AxillRp9SgSSlPLaC6Om1+vBOgKw20t+iPQ0W6
HaYSLk67UMITrK0sYg0wpJKXQHjHJgTYPF6OHMnjPx3DQm3H7/LVF6M0wk/B64T3
FWzyethMLRA0LNc10KU/4PR9Pge4lKHM/G4kzR6EoG8+BfIMSOgZnDadta6b9/+m
ZMdB5v2ED//e4Wq+UzcKH6MD65dCIxO/mt0kqutUhDUTHeKl00eWvAcA5qMo/ta5
OWoItVnFmCMHil2ydCUwehAmhMTtMNBmRJcv0nXIB8G1Aai+11IM/h8aSbXU1dUr
1U9NcqWo+8odtARbIxyzhLIqCDPBa182upCZkTdv4H7eGZPYOhLFL7vgytsOqLGs
iLB8pYesbal7J/nvH1AYQ9vYk+1qOcisbPDJKkZT4cX/Mj88U6nRwWZKRzYQH9NI
IwPhdtEuUI+PCDmGTv5BPs9cvfKUPXFLonJmjjh43W62FJprS+bqmGicewODQEdW
BqRAm6cR5i0QZ1DWxDttPciBVSRPn4Uf2WMh4xdqqTotBNoIpKO8HLseTy7nj7UH
5IlQdbtQnclget7FGixsWVs6AF1URikHdG3JsIf8UbaKK6TTw1R6WuqMtxTNcY+W
dDHOPL5hHjVv4IrlfZJ9RTMIyPbWAMo9/7XRR5SQNU5bS97kN/qlY7SKOQLOsW+R
/Ph3sfGJ9KS6uasbe7Yh7B2+7uK6P+eMs1Sg3tOoPiywIY83yCCZkt29TBMoKjRM
S3paNYecRk4NLx9F9CSc9yq1DPUEwxjSS4irmYVIFW8lHXuLzrHPbAFkXh1mqFZu
5a0c31X5UdQF0LuisFS3hx5v6GqEf33UzCeX5BLul2M+4Frv5WXU7VulZvNRy8Jl
q45OjVKWwL3COTd1kkeh/7Wzq3+8rjkIy+Gk6g/pbxR7U5QPzdQhnGNpBvwf1LX2
NAoPqO5ZH9nz19g/tRKg44FTdiIOZfAJYTFSm9PjILYfz0xn0+MO238cRzu1Z8Xt
OTPaWAcV1vvzC3YpspY2pX8Hf/046idyylDnd8BvLmhmrUPib2YSg2kQth5YphCz
MOSiXGKKmWooPQqM6cT4HK8kWJLYruA1pxKlaZd6FalByWAxlLr9UlSCZN/9DQM/
dquabpLJ7alFouHSYWmslUCl5r6sq+1036OBGh7Q8XANGScYPICfBQvqss/2irIc
vJEi4lKHsUUx7091L7qt/gN3XIHTghvCwyG/iUGCPxEdLWbWEEbdXwnPmKviBeDt
SeY4T1JHORE00R63FZX377sIweYtP3SozSvbxyzy7EiMfaNQSpb2J4wLO+EwJ9nR
ZUfwDfJS9miqi4lphQu89OYha7iTUFLVGFZ4dT5z0/Y8FuzKhZS9k63s8VkI0Py2
vzcEjg8Bg0jYyxGp8boP5O6YzuKbqvw+fPacTPgYLIs0sAjTLfuFBJ/rWhdlR6JJ
35PskqCipoOWbGd8+9D8N3m95rpxd/I3uKZ3DX6iSDFRZOytOilRBR5G6s5VReq1
K+uMA3SsmB8ggkyYUWJqqg8CAGykuTh+UxMAxD1HP2juMZqXXtCCtyHcewhWyr44
bmukMPosp5kSuguc63it8p6NHrho+uai1mUXUSFjJYZnkjcTxWVIBRTsyDTzlh9O
uwZcxc+YhYDyW5JefsYArmS03C3eYWl5AhzOqynfMpHBg1J850TSmGIbo96R0Kds
Yk3i4CHnEfG5jE/Bh6T08qGQ6AlzUlnavY/TvJHo4zTtNH5zy6NxgD3VK+nq5rpX
Z3Uu2vA2+jMaDm8kePqFB8hAW/+ek9QWRj6Ld7TCVecWd4SjPQ+8CCrraKDn0NEu
FKSu/5YH9dMUehkOkzk6yohldJc3q7BiM8bb92GHMy6SW4ANmBofsQL4OeC3QDQg
Cuf0PKe56M8Lqi4U8FFYTSYjvWlj3OuhUzMR9vAizVxOG5IF44wmUOq2CYTqhTBe
wPpa1ojjOOea7X3Uzjq4ZERh8B9UqonE4rqPNVCGBDAdezVzzCG7/SmgOptINOjE
HA4Djnik5T0vLIKKBAg+eaWsKR3zNl8c2I78sXnxGMbovV2hZzzhl4y5lWKs6ttc
oz/ctjQEKftFTiw4Q+j3UESAM8/QvGn+hC1r9mizLv19cucAmtVz/VUeyhkEzp/o
RSXjA1AyYe7kaVSWcXhYK87Ml8jr4uQVZoMZmsS3jhdroNQZcdXdN/N4TV5AlGhe
4/CNBjlmPzgVU446lPnjHlXQHjnc23euReXHYb085k6rG24O0NPJY0r5mMVJs5tF
MCBcO9HKKINXQSIQfanfmEt62pq1Kmvm9MOwxBkgJz0mH+0KKCc8zVh37Vj0Gogy
7YOjZRUQE3GzxRfKLIazDroOlMqJ8Iy4xi1mbehleXyIGXmewAmNsAFLmxFM3PbI
TYRh8kaWvTQIFXiPVlmpVi7/eyw6J4qccRDAoQkQJryPC3ljbX9eX5j72pBCepCD
/0NfFfUA5zoqcBYLcI1hn52kF1XHeRHNfYsLfWk2XWO6W37+XGK9khnc8A49MCZj
vHh/FMnFhSXfuimziD+Wc14fhWP485MkvqqCscsIaSH+7XZQqoejVI+tqhT0IGO7
wss9yZcKOqJEH5Ag/IBKIOHpSbqfprmXM1UdJPHeql9MCvzHwLjFqOnb1T3k6PIH
HeCqOq5I3lsfM1tVQZxVlaKtX3weQ/p6R5Do3BWTxxLqtOgEFgDMXEhN1S395C0p
IUz57kkod0uV9fbE2efyDcRqOHcTj6AGKDVMm2ya1HvQD8YksPZrRO2KgjKbJuBM
QvXlFy1I64sMmQR/gm5h+wI95XRjFI71WhnPTflxceAMH/Qa4St9ElGWwVbWkmgK
hrhWKOHgEqrNmTLWeaWi9lcD4U+QGGvvC5uspzbYEAzxP3oT/+eAxZRZyKY2nVJK
mAuWBYeft8Jqbv4yh2XkvZFEzFRfHALMI26p5pD2oHnX0jKceLI1xrXmCk0VX9cm
fgVoubzxd0s1w9ZLAmpgdhJm5Ng66wl2Aitmhkcrk1wHF1K51zPRwQhJ8E3+E0Ip
ZCgVmEmPK2ran9NGCY9InyRJ6nGZ6CdptmF5O9TCV1Z+CtR7DfSBq/mYdDMxhVsQ
aRK/RNTUz79DUSvM9Kuz06GJrwi4l5OxNy5ut+86URRqmGXrRVDYqhEibNDkej49
HBi6lGvT3+khJuJTaeg2Mm9xKahHrgeSEcjuu4ovsPVTMUQLO5QYra8uwiDP/Shd
EVWZsTygATaC5R/aIaorbnSDy3U0P+EQaCoXBK6J6e0KGKp4Rqc2Nx68ZDGxUBcY
1WYB9pVwyCpNDprRNAHV2/0ImlGCvMmoIElbeL1Dgi1gC5sYIpUvkyUApU/Cp8Pv
ZEdIV6eWmGXTTY8RW8GeHoBCAiusp6mVmDV+cUO0hXZl2OWIweHWk1bhd4wscaD1
V7RbQnFei7OscK78rY6ZqctbmjjBmjFV/Qi1sAR6SpljoDUV4dienWSlxS9hJzRi
6PDOeRgm7XDv02VkQL0UkMYv2T5SVkuDoJZlaGmLGWNQnvf1uX/Chiwkuw+TTKD3
Gmx54esuqHt5fX2Vj+hYEjbrZlBbeiDsxNEJxhdPJQjlIjnljy4R5JoDMF97VuFi
jmm3V8DFpsKPp0uVaHJ8p+01+fCKWCH71os9dNgSH2JuV2OnMKOgI62oaIFJUwB0
Wzkv2bKjwHGKq9Nprhfw8kSG163S4Mg5NuMonvimc4YfOzqtIDxl32H/Y330RYGt
+geaZCCy0CAots4QFhBs6HPO0oeGMFP91Rf5hUFNZCAK0OqxzLZ0ENQzEFzYiQf4
8uDHzAsWhyZ+VjFgmT7xOSzVkTsulQ6OnUGpoDP104scRw9GQMSebsFlEPZqOWZC
fsamRn+xn8gLTeYa2DXGiQXyngLnBaWxNydprUKtnPiDQC39fxHIVMilnFFePbL/
1yPE1lCyRrecljbegIyl2rxax0oxEosWhKbBbdtBYVIqYZm3UmpD7gedJSgi92tg
LUgVh9vm/X42theHWc04MNFuTPSsIQrm70QRmim1QTRNNHELIptpRF1v9LL4pQuk
XPdgSwnFSpmidJrXc7Nc4b9IIzd04eG9xmod+9pjiIIvN/EhxtYwd0Kx3GChGahI
y1fR4Gg0PfjQXhJrHy+YoV53qLtA1Aqo7hS1oRdDp6KqzK/gkDBlwqto6vOqDKAv
JvOf1IBEsKv88woP5X9VDSmzfTisbiLDg8jkZPnRD9lz8s8/Vury7ckkyJrWNUjC
pEvaU391OM8/+StQyJq/CMNrSJXgRHU6/Co6QtfmyrroBz7JMPbt8fjZQxFjAX8o
AnHcexaPbmCH9Vl6Umy0tjXy0/GETNmAI6+D8YImdLWoZCMt3avDirWujHHdW2lP
WSBFblaGczJG7YkVQtubBhao+Ijty/TE/XvcTn0OfxbpnyQX4t0bwEarXBp7KnA5
v4m3y6s/ZEpXNYh5/7vxDNb6TRlRfrZatoVRNvITPYL0agFKia4hVtip5HjgaIbS
pjAEtau6UMr76UZR0lPJkNQnNVSVBgTaF3mT9dCcbgP6YZmBePRwnq4ZO2XpE/UH
8CxO6pFltBhs1Bh0s7glee2fyLMEUSJV+BYbvA9OFYz+OrzIA00mf11j9xX/MtZO
9ysE76ysHQKjwTyBm577qbusyAID0MHurHs3W4jWxsQmeHEyuUq6gXLyXZx8m2BS
f93ucl3Kb8uz8ayLRezeXzgzG6Kk/NWQA9DL5k3+oY5BrRdz+Jjo7etwRb9h6ERh
FoZ772WG2DDUIzYCPj20hCnyT2IzIZr2cA++pgXe/ULi6GTPXL6OdrX+A1MtPDWJ
8Vubg8zPyzCvGpBgn4xTDUnQ2payIEqy4BIDICyehDMztz5EriQoP4AoAq8Eh3AT
MHyOwS3lrGrT3KUqqzo2lch84/tNSVK62KkdhWCEGfOZJvv8I74AbhuZzHsj6dmW
K1zFFKA6W9LthKpbAD4KbTpHTmuW6pZCj9ti5u9lOcX/4T1kD3j4YVeZz0S83xj/
uTni5GP44G17jR5oH8uhtJUFg7WyaKvmN1MqRk20OAinxbpkYHW8fCoFXgHB+R/2
+DHNTletQRetepYOMKH7w85ot6XElXFVJx1z99eqB+KwgnuiyUdIBV3sN26uNrFC
2sBzPf37/mN0THDhsK0/ozt+NyWF+vu5bTvUpZCChVi5ch/sSMlqfxuqaksTc3go
19K9HsjHePfP71zvDPESnfztfSfQm9VDLnpQS0oPr9dVmErx6asvEvc2RbuyFFS7
e2i/aYuyqp+A8Uy8Hialgl8ABoh2sq82KLCslYMmOq9TWfP/AeNb0cC7oERG8f0A
Qt8ATIDnKaJHa413qSjAVIs/CnA0w1kanqphSNCB8/EIO+k0BOvGGHN9xOn7liZ0
LHOWsntRegR2WPl5Dniga1aqz+P7Jxc5J8bbaPZbvG8I4RIr4+M9lud5MefIoL1Y
G0UJw457c0/bwUDzka2F7GCWExq9GzXc6rMRvcuxkbxhS3BY+SicjxJOO0gXbnka
4AOVnAneLtfOeX6P1ghH1vU3SJ/2sHJkTWsE9zHj/a/li4F5qqwtoRWG+YYJYiT0
SjSgFPLLcs7BII5nbE0Rwtw+WKEDJg9u2wt4vy6eUyGUV4j4ms/JSPoyGHLzIB9B
a9ZF6Eew0YbU0nbibV1xUHL/Qola8mWwE9UvRKmb6nQArX9PuygaTm9ipiqE3D6s
3kSadCjcipyg9P1KklLVLz9s6lx6TFqhHDl1O36UXucUmB5ikOVnAir7/CtfOkbD
HkO1jjp7DfyTZR+IWruylQ8asBoG9UAjZlKH61zZULQMsdG/sLbWP5CqRqx2+acl
VELw2p/62v7ZmR0VEVM1PPiGO8kpgPQ5Rs9WuxcRdvlBCdhtpRkJ5UFaO53TC67t
SiTgpUjvq5Mw4FAxIKDm+UliQJ71As+rtvVjuskwxYiG4Jegoz9TbpO90GDvxnGv
b4VFwBBRm3yPGmbKn4PY+2K2oMQXuID1nWxZ8sZfxt7M9OzLbDmIubMCuw3Gx2JU
E/H/yGh0CS9vUNF2kDpxGpuPZxP5ik4gmiLMCDBN60j8Zd87D2+pfYK/m/zFXwnj
mdSugEiM+i551W6cPtIZ8I71GD8d8jmyDDb0TEgymKUNz3pXzpZHCalXmFxRbd9T
8YS68LiwsOm0XjIQqCLQ+AJ2PpETecwpqQFDl8+vYHuM1a6dsmE3wWq4yeqOx1iz
sJaXz7atBz45wOLe9276m99DFJsRekRTR6+alhe2QIe2QqJwYwS2S7kuHjElnG45
Uo7B3cZuCvF01tm2dzJ3fyQL0q0sxK0Szr03XXrhq4Zn90FuzqyFPfuMJg4MLXzH
8gah8RKyzZxKiKDR+metvGgL/y7dDJOD01duIoC8GC34ueFOqPtk17ubm4JTLicj
rz+tAXrTGiecb7PbJcbnXl8X2W6qyR7jXxSgaXmKWxKI5dzhJ91DxfKBRhQL7xJL
n1fNInz2IEQxJMISpC+BzTjOT984hWlbnbrfGmvjBYT6NifVjgJNHiUwFU33kn/3
L8fsF6jNOZHNZvbTjTTmkY37Bb1dsFsbvCX6o/NbLrrockhVeUO9yRFtXgCd16Zr
V41EdL2C1hr05k387WLVS7FbMysID602QY0wzk/6Yedbu3J/WbhMpKe2jK6iuWBY
cJPQotvPb3rUgjKqZylxqanlnrHqIJntAhrUa8D8fF59nITRkxCohzjAWs4AlRd4
lfhvxM73FJFGzEDt2kVY8qAS28JYqLjwlyu3b8OtO9FdOUQ34llAHb2JqS0R5Bac
SyiK0RjgfCWIzW4rWpebxSgi+u5qoRts/onoeTaQ3hTZzr/Y5zD6tah9re7KR/nu
5bHGEX74fHwe1rI3/YnLcyLgXEzZTenHeM9o8EX3Xq53qeu9RZeqY9IChOzgSlhk
2ZO3wkAjV9NDXaYKWiepNw2Hi33Ny8InXDFd4aSpaUHyPjDVlZZJKRjKclUYsRBF
8/dvOYTlScBJ3H9m3sGWryKnrQBs2S4SIsavoRPvSu01TustW5eWHHhnszM/lV/k
uTyZrOUEWEIEndhhRjK02F/m95hyK+luH1CGOC4cBB6CdO4gBpIowtm91Wm+E4OC
myZwrItsI/3SP6GsQH0jq+5dm3GEKTeJ+EmfiNgtjtKkxGvOLsgxRnEn0MOhOKTl
NOpe6QgccgpC7zpzgpb6esVa04EWV0Ld+MKJCJZAALbAMGVtAgK+JJR69ZMOYOOG
d2gaiFGU3V01eGAK7TF9+Rd0aBqXbt8dDHO9fp3qlgWeVaiu/JvXiZgu2X32FCTn
Z2J7JL6sfbsAz+5ijgQu5+LACGje/FurH3r29IwrZgnlB5N9ELvC8z2Y3vBqBzkg
V6x9tM2NlAS548IVc0YokKiTxg9Aq2bUl/ok0v1lPZW4Swvzgt2OijgHxUxYSDwQ
5MurFIyLhyIT+g5JWXelupYoMXV6hMlIMfONhh7ZjdwPJUj9iAkE87Tg6AXpF0+h
OAvoNjbG/CPOqLwqt2VWteBL6egmnlqPVaZCuh+5MC4H/vqsgj52hFYrp9Ms6zaQ
VzN5K+atGQoiUltYxnow0oM6HyoAcTCxFIXCgrm8zk0l1nk45EXAm4vu07OE+T8O
1XGdkIn5CcIcjEp5rBB1/RMDZiIvbjlPs03a0yFaL0UBxCcXAPZDVK0NMy2DaJKZ
iIj5TG8nV66alLW+xlZXMEbmiNa+u6V+zKWV5zG8xD9OImRuIKcIwj7gaqVOQSFl
O5wZ/LfzAdWrJfqC+Ihjg/5PN069rbdSy0Z7Z0LkeNjI4nyMqxyJMrb5RdmKfI2B
p1Ct4ghHpAG3z+xrPlhEdOxlI+mr30Am45y+9xMZShuW916iUblK6a44OMbxgoGi
0bK/JR7nalji3f0lYVLAuWm9Pk4VyKmy2YIbEtiYWDgOqo7slg4APCrFloopn4uD
fWKEf/iEeDz44Mx7G4AFR7+zn9ahy9os3GYHLnGMxhzqbiu9Rq2GQv2801du8bOk
E0GRKlxfVESG5fDcACjpPtZG1SyWhEK0PnRt5bDzRIrUQSsoKNT7aFjvyIJyNmyf
bmtC25by2yeMqpGj9EGk6fhA1DxAiWxcRzzP0rpKVS849EW2KcLgvH1/r9pzDoa/
VFVyLSp4OC81SDCPU6LyoYvY8HJPam+1QOOEr3npOemnCR7LDETa49e7Ad2ko913
pHsnNqlYjHiW0EELTYpi0PmOpXkDP85ygueCd8/U38XXy0wEDmlkuTpZRsz0kDRM
ZUcazXsjFzj1YfkBPiaaATLIUNY059M2cK/ZKHidP2nW/GAkA1pEN5OGzpi3fYWy
50Y9zYtjs3ks5quC6OetaH+7cPavxOeJG/GpI5Y30oldm7oQSZ7fXfxWekdniKdK
a4NSgziwq6SmDfh7yGrn4tOogg5Ie2KX9N3kZDHrTJkgeACe/y60OA0aRFDsRtOh
bfisFHh28jbByBEgqfHZUBmX5GDzjH0WAyMtzxtfKfSkehdazo33NsM+10O9GYgX
dDjb03vRHxWsfb2Hefrh1AeP0e4Vr5cl9PAdh0XZDVrXd3g/ZV7yZG0qTEiC3V/K
c53+zjJp8t5QzGCBUMyOzFS2W3d6kNx2RdbR2wT+JvfDqkii+ycziwRgwL00VTSc
LqoMqFqRjIHPKwoIg87TkDGkZ7NzqzmidiyZ+cdKT7N/T2CJFqi7rYrDIm9ndD1Y
TpkOSQ6Dndu6MkwwlHc9WM8ADbP5MxZbtrPHUTMujvOqA4idAxwXrG88wVJWEIBe
6PbSUyAsr1lqi1HgfCu89zzMQFsti/2A2HG4gkkO0JNVzKhubtfVK+s/BR0xbGKB
lvYqqEjtNzMgW3RPKMS8qSLV9vgh2bWfdfIDXtIVIdel9X41JeqeQ9LwIQ4oPjcP
S4v/9b4GMdjEcevbuuTWByHM35RkSv+Yc9VNb1YIuEvkKZSBQvLvzLvAT3SWl1XA
2x8nMdjhx4srROR0pw37dJkM4/5F7hx7qeYlnJf2dC6kL8JSkTFGVr7yFuBnzI+J
g3Yn2zAapao8oYIHDK3refk0jlnrSmnZQWj8HTZvXgeUHZQKyfwxZAVZx6E/Q6FZ
O0t2DaVeTTTL6l7u1O5UoeDPmsCMDBN85fFV2J4MJZnYmGe2ftACeGHgNqZad+ht
fU3N60gcLZhg80/NIu5i4UF1pnBNZzsmlIGS5Xsg1bwFWmuRGqdDaCA7ycfbvIOl
efuhnUT1nTX1hU4IoDQGVUvhT4e3LVIqIEBdtRiiUfiFHozcl+YZFGucFmcW4V7p
Sb6s4QZPARtqK8rAEoOyDtPHxEKwQ+F6Alw/X74/61IyTzV7tM67Uj1ne0o2Q9DI
s1qFFM8Cutfga9nSF/w5atym2cNIMMfQXDs1sMuujIc/kS5M0Q/6+bYE+Vqwf9M2
XtYS9W5PJiTLyT/LYT5PWSU0CS0lO0WzIQpYVGXVUgyqgCD1qK86HR7Ko7tCQ53Q
Sie+mYCGfHhNciOYFyYOIGzo4e4u6QxPItTPGrSVi0YsUULi1s1T4xkWSB/7VVn5
mcC6qwlCsSYqz1Z2Uhqzsx94cyCOxwE4rYeCeJ4pvcv52jAxA0i6NM9imDZlKv8O
7tw/iBN0CywURf5nHJM/6wkJQ16Pw18l4/SGQcY10QfFIX83uDSw1lQtU2XAL0mo
G0cPsADyjgR+NJ7oa6ZHOKazzDOJXVnDGIcu6BbAlPeG5anFsMqkPGqlhE20Ofa3
RiftQqGsOaz3i8XI972t0kmQ6dSjBBkS7gIrio+qgCrU+fXbriREiRbyZ8jpCx63
dHD1mAAgqcOkPCVc1El7nQE7HPbvsRU0SrCBelSYECGURI4b7ZZwDmiCTJCE7SIn
aTrQZSM3anqijp5Us7iWe3kOS2yMTjyhuno0I7L2IhNwLkUtg8sIFuU31Uy7Sqdi
vNua+1CWxecEojq+W3tQjbABP4nM++bdhQtCGfD7JxzLYcgVD4BW9GlaayFCQk+U
0OAeVCJE5rj6Qxk+d4uNmrbQjxg4vWzuZQwBJ7OPXYVL6LxjSwvLBlQubXG9IsFP
edme53NOQfsSgZnCs5yqWB0/hk4WnPNe44D5NC29xfJaeVtJth8MkpAtjbvRTTb+
obXai5hLAXEhcZ3eTsMdjGDfIBOPBDBUxwXw0VqbgZ3V2HkSTBacdfcTS9SzVQgq
9/ywp0mplUtan0rA+X/iBfGbTL1wwCL2DqWvVa9wGLf7FfNv/9Z2+BTSO1pO28u+
GgxgPixUKKG/rBoOkX//f5Di+EGPqHKQNawKsCo3pbU3k+gZgiIIdpHvx1Qo/zVK
1St4MyWcWNfTzcokHWvNOcMq2UkAE+5lVEpjDdK4pn07r6PLeTc/Dcu7eRChAjW8
j1UGRkUzV1O3mkpaoxUyN0/1+lxUw3RYt+rrS0QUSBkZO1b37R2dkJQzbem7Sp6D
DfZNbefTlvePPnzgSPaoirSpSkwY9lZ/ZA4seqNPcCTpQAWZ9aK+qf98njhfddfN
KJSAdTUOYHX6wRdJS4CigTu02I4kQwhZC3oe2sjS7D18g5urrqGXfXZOvf9zPv97
bi6+uJH+g+YuPLTJN3/UmeuFXtF6OAONzMzR/DYyjAV2LNz+IsXX+jxJwgl9jdxa
NcalHMCyLAmMtV1ulW5MHix03W7si8ZhiGzU/+pNYOx4T63DfnznrTX8ZwIZfJ6w
BoUb0IqJqYPkdG56FBW0UYIqTekee6s4q+amBfS+F1614LEgS0WPGKQXlkdUqCJT
3BqYRs2/UOvSQ41J15LH0Bim4IM/l/61HVqRHJ9DF8oPbzy3KvuhKoYcxgl1UO92
tnUn/nPqQdLyCYpGJZUhMDXkbxuXTaOzCdCk/0bbIiz+hqaNCXqttN2Qu3dIGsja
uyT7brxpmtdnJ2pfqj1/SCB8ZkPteYbBhGroTWdyKtRgWMC8TKEABBEgH+01iSgY
vfGB0AL9KKlJOhsToe8aXuI7M0LLfXdYG7mHDiHrux+hea4Tbzy+JhKiQsxKpWgF
jxdmyrNfN3xtYtUR5N+3nTYN61ShSgnebxKuOu+AlKQo6KJ6X2c5UhkY7A/wmzkF
plsovD9lSLskmUg3grz2e7UE6b4rmTlYmi8H0HhYwt9MiD7LGEc23Q5n57J+/hW5
Lbd9R0qzj77jDycY3nEDz9hDK+GtbzOEzkKyZUd3/rJoJoHSnJlGiucexKUlrxxd
lf3bd0LEMz1nURUdJjlQsquk4lXU6kKZyq+Icu0Vg7O4j8Gq/77Ko1E+jZt0mNMK
fgyiPo25ysvTpmkKjOUZrSW6/EdCqNfgKDLsDfRODvTbQ3r2aJPDNqyy9UQgBfwU
I1+W6x0nmIWghrhKR9nG5p65LMor+jSXFWJt2uU01IA2bNkZEvO0/8yAl9/g0aUB
9xKmEZzxzOAGiU/9WCmGOq9y1auK6Aww1Gn5u7z6UwkQHxmOfhyD9nWGt0vBLy9m
vTv1dNWzGrziSrSNJbmCX8WNnoRBUsXcA2UW9vBnNWUpP4xY+qNvG6lRvbtWiqAQ
tnoUJQXSpCQhvdZVk7agpFsmd2v63XZPAPv1fUZAD7SVKYaqTY6rqioemmR65A2E
6kKGoZSvuqlwrqWBiAsHkp0i/1wFB9MLe2jpd577+PBVyqeY6FPRNPa0bxP5kpxr
xibjr1DN6IsiFZvmfaPRCf0C53H2MpVVc7AAC9cK+Mj9KBtH6BmMFBMG4RVPjhFF
oCYEx0gmVKki/R/Xru0cxtLVAlWs4jtFPmCPowWb9ycTcSwscrLoAl/UcT/iTo5q
oToUkbpcguFy0fvXXVT3+S6fufJ3o7czMSUJyvfL/mke20l6ex3U1PeTPE2x5vTL
58us7JEy7kzOnkEU8dxhT5v3o6czLVaxU+p4Pk3svS4yJX/o9e5V/2NxJhRvLER7
cQRO8fBYbYuXqmB2igHU0A/zJLqshxrHI4H6Ozr1nCGcwVMA2LeUhsTlPVpAjdgY
wfvnuf781SOIUUjkN4v9x7zCGnnxhctm2J5+Hjq1sZTGhmjSbLaLeH1SK3UnroA8
lNXw4U69QbtfQYqWQKrYqjPDgK/C3Gj9pwj4J2+E64mRhOcPr+6kTo+h6CXR3Lbj
VIr7X4xm8u6Z8hHtrr2LaPUZm+0+ZwHS9C82lXJq7+Q6qHmyo2NKJ4x8mDynsdBx
6WHtX9pzbHV1Me08n6AcjixD9u324dhwPzuNIrPpbFBhMmQGXjIW0Tf+rxgZy9SX
zIegLwfcXcqkKbUc05TMfxuCX+cUJ4x+WN3EGTivNIJbfgr9dTn3TNlv52ihONNA
V0umTkcFicrqjWT8/JQgoMlt3q4+gNIsff7j3yENMs8XXGL4A/PqdkL3QhmkBlAx
r2c8ebvz8ROnmjnJb/um/wOcWkNpP9muFyjAezdlR0msYQT57+wMKEAJD8xAvH+G
deOrAJxLRLFWTnNs6BvbCexmQIMdAbyAKuIjMDXSepvAtw8YHx82EXL+g9meVN42
HEpw7/SMYS0CExxvpW/Ypg4HSE+gPjsSq6+SJ3g83KO0/H8QAJll+Uv2zGj0RXq/
zJRkHDEp6YXWUG34q9EZXfKiZB+SlZfy9Po++lZhM41qU20zMF0jDFlzRmaAB88r
7YPZWXX+tXzm/82ZwG19L2CR6JZ2Ul2dexn3S5wRNJSr2oXEmHqUUx9chh0Q5PSS
Q3lXsQOq3+UYBELEPdoB5Oq1OHXraaOxH5QnlQa9ugaHnh439NN6GPxxJIpJFhXl
avBTpS5o/MrYzR09D2O1QtKGUpnSuJIrRJ/p0BcL+RzTeJWF3sfRT0h9yAnTr03j
nTYPP9IjTkuexXGrLOOJjVO7IQDsHDChFVTsKzN50F/rQhXgR4PfK2+M4ikJAKx7
hzHWY1JMwESFocIZLls3+df9hTEeOc5lxsKlO0fUnonW1AB/53kNDpXuscbkjunl
buq+9EyT+Q4VIajxqsTCydWkZiwMj/Ek0Iwalu+NbV1GuOcCc5rXcG4kX8qWefh1
RZSumKLzA5UoeZBT9+IvnD6CkGbEcud0jJCeZdc3LPs93Dlf6Jxpdt+oOzQFC6Jo
Kh1pHJN22UjyxcfJVjTx0dQnH2oHzuAvSLE0O09qHu9fFYoNvUrm9hsZKtbESSNV
u7N2gzDhS2/6T7zDHpRXk3wsPedc2b8yU3k/m84vdYccWUt8DYBrQw2RDioLrgI8
O+zxqq+FJYEF4mS4MVcqZ566AieBAsgh2XzvqJ5TJVkHJcG0kzr1PwlI1nRDxBPr
6x9P9W0kQmm93gtQjQX5TmpcLvVpxHTe+iOxcJsIlTqsCXgFK2jYkftipCxzg1BY
/HHV++qcP/Ma+jTWnWTJBIn9AHWkKotXGQ9tcIiSxbEXdR+6ukOP7IsQsqMcMntE
w7n7VPDl7d8nwKpPbP3cQgDnEZjlhG6bnTam9S2vufEKwYWqd59+DXo2kRnnCvXB
loiTJBfoYsNivO3YQxEJZefsnqevc1+6c8J6z6jR53BEpdOCAPI8z3ajJJFfhfRN
O9Fy0Yg2mHNUL0PG4YfsBRVjRiUx1FIs0yIfWEpuNWx4n6/XkNAtrOUOli7au6DG
IzaqaT3Eha6Vjlg9rRyvHjX0tcg75NOGZA5CUEqikz2bt83yzsF70gBvW7fhRKXi
Qt6zUnPK+9p+8KGHwWynKWlV9T6iuhXRASfeSP14vZ7326B/b1ROVtI8Mbg97b37
UnQg0wf3ghBtf+ydF23YlfLz/0uYVS6at0aTd7sz9edFbP6rcGIw4yE+dNdQux2f
tjlmUu5bXVCzjF0N7wW/dApzMG11QZ74p7Ztb9P1FERvvR5Zok5GN7svZIQs4pQp
H8o5acTVl/RJABddAKyeNjfMGJg3XbAXt9na28IKhGxSHRrNaZezq5HMRGc6jQkc
QR7N55x4EIc1VaZJv2dV1bC91jmJkek95RIKIBdBX6FDORIQE4Of3weOgMns3nrb
wbm/qzxHaqLtk0qWYa4ThbPGQLX3hd/fCR/cDxnzbayf7bhmLTvLPgowPiGAja3S
qvYCWyoVCqngWxggCqMHZylkeiYMExoBD27TpUbqG+VXLHWf26BI9BOmL77HX2qY
LqkYXmUNy+6pWAIxB1sCT8G60wP0/QwG9AWiJ8CHBoUY+JdYDv06wt1p9g1kspmK
6cO+f8mpzuXwFdpqKxGbn2w8lQk75YpcuEcrBwUQKJjWSLpnduOnVGI/h1slmwSA
VxTnOa8kwUKHsyI5TO8J2yjH5NdM2gJkXxa6OfESusxf7HxC5w5Vu8yqLehb3hlF
75SDWGUSQibuWhGtdQfCZcmeUBCwpUBAb+Vjk9g0pWvu2angGsgZAmrjplLsrFtq
nGhu6ZXA9P/9/ohHrmvheYgUgyp3CLgPqxImJKrKfWqvvsDRXKT9oaEbTIx55Rp6
trMVDZ2uBH60m0+zxajr4nwgdBSsul1o5dAdi0K4pkitietj7MdQipJckG+7dHyD
dM9/hFzbESw7HjinIqv7WCcYdZu4rDIJMJlG5IfPU+Li/NwVthMTztsNa4sHnYxG
B2Ll434Wz9lj3ARK93O9O0iFVi1D9WCP0zGCra4q4qHGHNgKSWHCk7bglUCW7Dc4
EfO1aCy791neJxnMWJRNfavIqzrwXUcPSRZV0UyTCkqzboGKX2SPGBDe7L4N5T7w
aeVlcbZBZdJkPhSYdJEQfQ8OcWhoy3JTJNvu7Gk+30PUZ4D6INIf3MJNUc6/efD1
fl6K8FQdBppMS5X09pScOy4gUi3hFq62eVkhytuOsP1Wgm9ct+uwa3f3kCD5dvl2
h1AVUEI2fvuE2PlN2QRxupjiP/T6n3qt7I8qbpCoDyIgQhettxmjAYcH1WuN0SXF
u7SGk4bCWMKHoypygnBaUtejNmv6VlQcctDiFfUkSmuoo+IBNnP0pq5v09tQo2gN
q/2Ewkh/8K6r+d9dPIa8GbKnSUfr5F2TgrtWe0H9+CdSYKIv9/R1yKkEWGYd4oP6
F7UYg5fE+T9fJcUbFcdzhdbxY360N1oZ5kEjLneLc8ieDrtItH5KEB4Hc+vc27D5
fQaHKVdHfRLDc0By5cxLn0fkI8EdB39P+rdT3qvr24e22jWDaQ74MjJoIZG7q3ru
viI6Cj0dez249C8RPNUffUNkDMFH5YuXxsz2TYY5SonRd0O6PsHbJQj2Mf08nFiy
y47VdR3CbPMfhpduWQGhrSCH8l4brFqnLQkgjwyfteQM7FI4ev9CMqC0/F1LeOSZ
0Oxtm4cxsre/4k1yAj2Hza3uOj32x434et8pF88jNDJIr76TRmvVy2LYon3XtIJh
Z6Y4xSya9QGe6r/eypotc4CY9uuTTjZRe2z77wotK1RgCmQBZVGf8e7my7rHkl4a
pNSyZIjcZ3q9D7mYxtPXXAOCtaJCFMhyfBa4oAx5CAU5Ft74Q40FKufpi881hs3S
n8Vl6XEnKVv1fuqTkCh1Hkk+j/pIsNQ3orO7dYxNuvxpUf4W/gWhzTS9LEcRsoTA
eEfefd797B9tUuFZYcdDnfO3q7Wc6aDTVctG96GvlafmaYLvOMnMocDk4G6TbV5w
dlAe6t8tnwnLUaUrLRqP62VkVfrrmGw3IErMrOdq0v2QvuupxfhKJW5ePojmAJ+x
lWhd3JGIUjcAlqTuBbDYNmM5WF1Ht4hGRAo3zWDtCP5R3jkW+8IQWRE6t6ba5L+k
7oQxqTJC86tuvuGZ3FKNFHN3aSZni6X5RgwCYK0vy9zrta26/NZPOw0qNzT9MyuF
buGcUZ0zKrr77naNnJdj+tdINgTkZLNTz5+7qG98GSJ8N96kc89dNRAwidkSwa6Y
zceivL+8w4pG6E+Rt1mJrAwgaifEfJPUjdVCO9S3GHbCL4zgWC3yoaKMUc/keMS6
4iGx2UO7XgP9Cas8kOXMll7dex51SVdbjfF8b1Bo6u4Tvqc1t2TSqSXzkQGnzdL2
EmxSoZ88hGVhBZ4q99SmHkpNvN5aAxCB6o+C97nCoDgR9cDG4qQvav+AmjFXORer
tlTHeG4pNQHeWpcoXOav5Dt6uVSxz9mHtXPrYUSjt5AQ9pkyb0/synyi6yrp6CTm
gqBk+NIVrtI+fr9FFD1iVvxWBr8SSbfWUFd+IZ4+ooUy0XFTllHCvnVbya98lC8a
fobuPQWmSdxWswzOKookaBEWFd/dDJmnvlzz7NWP6p89GeGXcWvFpqR+Ih279oDI
Qpts0EUPFUGGvw6MqgCZhGEWiHliTFvtapzQl8s/W51PknBTBG8xieJu97v0enlB
9cSN0uZ8dKsSgrY2n+qsf3J9hFT5KJeeA45984P5XsADjZUASW/k5Bs7Hw4+3k2N
PTYKxMr28UKXk3ejymxZ0eizSygpAZJvsWIqxld6uhyLJl79hOeVsOv+dByq3x6+
fQvs1oyUGepQPTyHYpIrGjcyYMK4SaHKRDGkOnVvyWJh2XF0vAff8pzfWROOBprU
hcMDHsxbjXkikMkbbGAzoiTl3Cx0/DmNRF1AOYx5ZCEvyTFixNGcZJQTnzRhGK0P
JQfAjwMs7U8v3BUo9XUAEqFq6QN2AzCWkt8/FCpj29SuynVosyrH9BnjECUOp/Be
eXKqhrFkfc1y7IxN7xjqKxWqXNZYq2AjMY+51g7Ysl3xHYvX9P2jKRcaLTl7nfuR
U/NdEKvoUNUU/NIcUVGpn/Pc5mYCSihjm2GDGdspLw01JWIFHfHjCYgPGR4jtcUk
wDpArFiG7GGCUNey++M0w+vzcWlW1lcwO1+/J+fFzIVZwjgAusRisSyQgxD2IFdn
4tpo7zHUxv/kcVNukbGZcRfXh9NynQV0Hjz6fveA17AcE7Q0axKIdtqiZ9DSmTvm
tEulj9X/7T/G47Af01IcfbRXkJHkUxqiiAUGM+4LhDB/Zc2sKexWr8V2RxkyaDVC
ycZhyWmNJrLxUC7S+Bq4b5yeSzZw4LhftEZvC8xGKp+yN6AI0DrUYJbeSiHbmLXU
UyKuR0s7irbxZKsb3BGYUan35cddZErpphxyLHg3Soh1cDgQWMww2nApnIWy8o0o
yZhHMyDqx10P/9qttuw+BNTfMsEh9R19E62bF+sR4HvhJzyjq5VOMK5PzVoOSOi1
UfzIbfxewu0x1CO1bh3EDTYCJf6+UrEgZu1Qzooc7TphXTqls1HCTn5D+7x+QMtl
yMzpBRHLUwRK0ui0owss2ljPLKKXsIdegy5+NxCeiwev4zmI5kwl1iDawoRyQUou
Qf5R/hReO60gHESZKohhWFr5g2khlwTp2+orRIAYz9nXDazBhKeBkjtpqSH4AcDp
jaQIjNuz3mILth/AqN7O4Ov+HFku3pGHKhvM33+dwjUKzMvGckvfSbr3wBeFid3m
c18ZpgttwtTCb7lEPxJuAHq/BaY3IsmSsk3bP/C3+osiaI7Z/6UvXpUBd6nDgeVk
JniVLqm8SmfSrX5pfa3Jens85QGzoBBHls7/YZEteenR6/Q/1UdOibJlO66MMR7w
MwGmAkSmGSQKaPiUZNopMKcaAdTvl6JQKqY1HySlVOqOAKJnaG1hl4LvXWnpjaU4
VQnllNC29Je7VJNNC6yc5x0OoWqkowYKlaCOmzeHdFj+8gMI+juZuqSPvKd3BJ+Z
Hr1XsaraTwr2SB9P0XDGlaEp6BgvFlUyq6FOckPthtIOPJojoBEUdOBGstGne2KA
/Kz3Y05SGjel+ytn+RLNjiNrqmZf5CsWPRUSGt5YFZ3lRgLNYkqts5CgD3+xH8qm
0y37okLxelF6adMX+7MwvWqIt3vxoRPj2mwQlMNTjnyG9HsY7VV+xcY3EF+Dn4P7
abVZrEOzZec7SZKEAw8U2oODfRWqqjXFnB0Efm7Vyf6F84entpC9+/LaQj+P3+hb
kSefYDnL88feCchVFXqv5byfCHprpvGkMGpq/sh4dcLEfEpzrZOzro/Jr+IY3kZG
hyo+nFSuvYlrsvlWHyIphnsexnpJr0g+biysx78xtpkCC6yiCgE03ct96GlTBXm1
C6GgLcC3NkM9LaTrDtGQaj4sRqPKaT529sBPrjM3hXPo1vE1H9LdEve+V9Fr59mt
//cif1f0EeJm+y7r5JC1Y6RyXmQvWrTmKCG6GeVGDktZYE79H96jZXt2JnZac+7x
5rH2n4ne2aaFooBy14GxE7cypleMp81DKDbPeNdFK7ieDBb+po3658OtzP5HVqWR
JPhVEuWUzZsvsMJG5HCBG/H9UXR45UNc6nGOmPbXKNGIKBJJSXj2LZdqM5fH1Ocd
TyttTTAz59+0frpBIBkICRAs2gaYSmLUAkelNSOe5mpEwR4KTHW3mOMLLtKAnKoA
wfCwthOtPEce1UoyF1p5mG+3hV0pqBJuSD0yGH2BCW1pKFFY8Ct1lBelpQnMCfH3
jUFyr5KoLAUOrL7eDynZ+NUMe4hP1qiOZOdK/9JGt2HGibTNOKGboy2B4+QngUpd
fDITkGrO/ZLZ1SmdWLbXggfH3LxppiAZZOK8GYmSrBSeJ05JAqTn0L7DMz+5IxWf
s/XQaacpdAV7mbAPVC8xX9FFAncpZ0skMmlHjD/w3Rtxn2w5X/3wI/Lj+2HPx2Hg
PjEL7PUN9Q9YAJNDtjmEA5hMvfWYia0CI8FS06TfubjqSwCZkgq/h3JlJAkEbZhx
fUdO2OvG5uAs82hgn6DRnPeE55TIhSAbpiKGN4MLa2WcRXC0oie/gGqNkqVkEk7k
oWI0ThcQywbfrPUeXEZHt3WHxnF6DJoiUp47k2QmPOU+Mjk9/HesBzR95HeS8gfk
u2qJ/qMlS/xAhdyjCXICLY77eG2YjiWiFC4MvxX/sTGchqUrrP9jN3sbye8DMRX3
ayIg0xwMmTKi5RsPodC3lnLnrB4AClkHrwk+scDe5OzQSCKYZnkdRfWVpE0fvNMy
28PZW62+njdAThIzaJxf8iKSqhzIJ+8xZlF125HYfx1ubczPtWtjx3HXrdtE/AYM
sYYL1knQSd72P+fmf57lC8Jw76vmHsZR7w3RhLBf62d7wPLiJL9Kh66jPy0jiUj9
RlRZS5fgoaJjC/9Z3XXCWrZq+1/nUrOS39pqaX8EZ/iho/LaIEMkrfMyYeuPPdjP
LwrTVvjdgkdzstA2NDL1GEny0T+rCpvU7bdXY5kYPqzs1FIlNnERbED6Ct0RxLqi
eEzodfeRo53RAu0uxVH7cfwuGqIIiTE2onycdwZ4MMf2LeX4hGS4PCiHC4g9VpRO
s0PCylWhtqHzsjyU/ZKP4F8wtC5CrJx2FIZ/gOgWTfMY9B4G1QIw3/RN88EgUscZ
nBqE3JJMEjhIEE+Yk93PM6zdX/5SsjXNiOUgpFEteoSG3gHFFn79n9qGDoCmYytU
pYqdA584FUQ9UuILNFqAIQytMfpzTayfN1OAba1u8z6jviXwKSGkIc/AwcK+2bY3
LlOzXnlZpbsv0Zs6zvzwe+2nNbFM2NvlBSFp4QTHi2WMJr6bKADdnmjIF8Skm9ER
xpuuMdectGlQvagVE4Qp8K09e2iixbOGzUep7CPssI+eOKB15l4Kgk213GJSptQM
JH/Djyq4pXCsdwsjVuYu7Rrw6cbiHtx3yUkrruQctOpYY0Pi2SY8NKuY+Xk66IJA
/FLx2U0pYz8EwkKSqx9M8qak4QlXyriGWJRPEjWzzQ4FlZJmoYyVDU1VN/Dt/W2p
qQcAsnlBPCzYmqlHT3HQkEylw7DVOrXWbMbFrHvwtBUw1h+EvPM6yGsDI7oIscsW
QcbHQY3Q38DQjoG+q4pl6rjqQX+gLkunZtERhJUxBKKx0K7EaPwXzaOwBeNa+Hha
eW9ypZDQyQJ1aZ5o0aD2cOz0lBRw9CrVrc83ShOWvlfQv9TSsGTpw8S6ImkcnXum
jRCuTyEta012IzREjPu1AN27cGQjOKhp+TLGJnyj0vo4r5Wjh5H21RFhe7WkwZHL
or6NuOr9ahVMkkEKU63+YZC7XxGWRxiYxD+WCmjTsgimTBAlgzTnJ7FETA0hldFI
DpUyMGOsBMR6MXCUOb+Gf9RqMyaS9Cck003Zzf/aNIDp/j5XXLCJyKGoPFvvcEdC
Fyne7ahgWRlB7MEAxaVWDhzTyvxbDDcZSS5VxxSEUE824q7K2ngjVkIvs/xdflEH
Cb9CYNsgFLDuhz+NKSUXUaqUwdHUBhnQcBirQap58S58dmknHzc0/4voniOM/Avg
varKY/Cq1MO1g5xMZYi6ec+EroJhAQR5RNZHglcYrzmVqw07r7GQ/Qna6VAKQz4q
OU5XD7LEcbFL55snbE6AhJWPI1bgk0iTF6nX8j8DdxOxJEqbh4IWO/SxwQODbTQ8
jjawGjFXV/XRFDSzqnLtNk/xrzwV5D+upJB0P6Jvwmto8Xq59t9sWfxsVeMp4lfX
3sLs4GgglRb0JqfI5A8vSROq4FRjQ0NGSS14HkGGZ02brP7aTbnZbWHlleu7gGR9
bKiO3AejVI7Q+jmvjbn+dOlB0jweZtQKV5WixcynItt1NuotNI03twxqEuAzJx0V
20uyx32K2iVCV75/Idp3P0nQ8ICYaNM6wlBI8mtBxe8gp2R2StJ+fdqrMXNBt33z
snx/yhGJ1Y8R3LJNRqzKplSzx8xmPa6+YYq9wC1IlraYa+2Jc+fuIBjHw+ske3/R
5ACP94epUDba5iQLiGf2yRVYDbbDr8zMA2xfT8j9kJWnAcde5I6C7thzkEd0Rc6e
oMRUF+w+kmejbmNoLMGnIJrilIg8Whu0c6VFLGj7HAwr4bdjjE+RUmVFXHHAHoDK
32Hp3fivPUEf1tt6i7IvkvZoarTd55yXagoAZuNLO2shd9krJoQOdBZFIKKUjoXq
d6DLoVmxMbwgod/0sS6Kyr5dSkF7lAqC7Bi1mZ67VjCdqCzdoxgWaNpFdNAazx+B
RO6HzjErHzusbZsOkdOFhjQDIwPSDNTDNdM5Qqa4r9wB3mqjZd+ZBbO+Ii0ADOV7
xTlVFBq5P3vIkrAu2OTIXU+ssRHqHdMEhFJI9PY1cr6oZm1fomYPZMETQfee8Ejj
xbqmLIqI9UmiQZbqBnMp0EmJaHxvBNvK7QBkcZXXpJqKpaj+E8Si2dqt7aatb5mQ
F5BDgW/QPkAqMEi4YTyT09fY1G2sZm/6P8J90EEi70gDjCiI3d/DFt9HiJP6irAX
Pqc+MIeLggGqMN2R1s6yvbppqSxBOW2VIOwZCd8vfYDscns+3H/wr04q2WS1jVlj
SqPCzH9AfpROvZocNEb2qGvL96/25UVu/j+hbmlFcY/U2tsfPNczuh+VALewVHJF
wXie9WQPqpyBAy6cf381RKXNyfGdEX1sHzq/C7n8XcWXmCXsf/rviE/mPS4uMpSG
wqxv/tYo+6C5LKtoJprdiHkuKX3los3jAPT/HxPHx4Go3+DJlKHHF5N05EFJ65as
TpwCPoFjAMsFyrgrnBmNsDdsUurV1qTiB/WdUqi52IdNtk2lsnhnE0jLNfnFsY3E
KYxqvG3LgjhWKIyXFL6aWuulXbK1UmoMiY7BV2OZ1Rmh7jhFUsRtX2lI+vw/ffCK
OBuz5Q7dxxJek4zLBsD6X9QFxNFaIQOWlfi/FoVFJn+vNz+3D9J8iV3r+v/5g1dB
k5ROrKZkOM4+le1GHjSlLoL+qynWzPMQy+pBIyJaNlDaUMIl74AdmtDQwbHGACX+
wK//aOqnGqZQk02KmcKDwrWHQ6kcabz5YHPAON3y6owycoKhEGDr+f8gLJOlcclj
Sfq/dN8BvMZnR9OQxsf6QRuVVUePhZvV6zS6rWCQC+Gh0hE4BOVZOJe4rUc3Va26
fEqV728paw4Bw6yBtStEF+bg6ktSfGva0qZp6pxEd92JU6s07ragQxN47FyBJ9iw
W51RLvEJMCiUxvprhHDf+lPbR0Mcl/l0u7K4wSDMSL5gr8hYok0+WdYI6c2T0pLM
iS9nobF/m4KEX6Yek33qkasaZHrgORnfgMOOcwUPHVQxhH0Iw0TPvc+9XlDsUlS0
udZ5Qosvq9NBMZDfwwUJ2HXOR1vUqENAmRwaQJky0HqMVTgH+VlJKVk7YtY6clxR
0fShUQ9re6n2L3J2r9t+9JwimbW9HcD1EdToPY1iqA/kMBorYoRI1qQ3u/Xif9va
z0/AYGG1YhMrjhXHzEafP/4UoB/20J29XAj6bMTVdBPnfuaJacqbPZ8MXJqHJaJp
OS9NNWVHBxQcwSN41Vq/FgS2tuouawtk5YvXX5fMdcBqOW5zPlO0hnQwyflcKFdE
3DGbv2NXbAdqbXye0N530V6KVYYDFqzsiSgGwmgmVUtc5UqVWVOSxYpoakVATEii
ygkzW0qjbbCeVzgXbo2Wwsgpn9Vz010fI00GBOJ0do9hlIkXBHsoO4Wyah29YhSJ
xKiXp6lb/Hui7be7nZxRZrRaM8SBdyJ2oUzKtZmkVEZs+yUFjrQdFZ1XpeYUBa8W
EnwNhzn6I3b6Feyii4lD9cTHt8zJIFgmS2h7WK8U0pBuUOxNwQurHEwhf4fRmL6q
9pnsZdYiEwleRebApzJFyFFWjszJuva/KdAoQSqv+e40CVcOlIBgz4PTTaGMn/H8
CfcoCl2zgvhpmvW/V6p3b96QavQcFK/dbmYDVqB2j2XPN4cGy4SpeEMJ+9DuqIVg
3im4EfVNfU0LbOazl6a+0PaMP1W9qU/ljvlDFMQLdsc3ee3ICioX4HdLImNsR9u5
LlINGop38UKH5OMwaDZnK53DdoPsEEHPsFNKOw+TMhIlwWWIAIGdcqWsPt+6r1Ij
+wb6WyHUFFt9ZSixxI500FxhFV8UJ6XJoOfBCW1vcS1PqNppDssKXHHtcZ+jBsAw
C2U2F97ItSZYLRQFJKWLFn46QYx5hTxXIdUXbNbm0UyY/r8eCBiNyIHHlIBx5F9u
UPhcuYw1AFjZztAEThmYdaIdJZNqcOoHRLCh3nlnU2+KC89plQusN5pKSaMTQV5J
9IDSVtFAmiojWQKIhGBiKRIZwuTcvXQJXHG48Mauzxsh/KM4fBbl4T2Ry8rEV+6Z
p7uzSQUyBD8OILRMNoUwH1x1aj7GtK5osoV5F6AJn7CEHeoifhEKb2uU3vdhsKte
F/dKaxvD+cmOiG4UZ2mHOVMnvU/2RKFKF+cTpsJYg/n2hTkIkxLCZKybH09Lvt54
0GfCZWARpqgGRLMMkmuShCN57TQB0zs9ORST12NdS04L4ehFbxUPlN/3yb9ReW8/
c+3Epou9o2DI1j+MfpIU03lVhVjIgWVcbYroil/3VGf6G6e/nCbLbjOOt0Or2r+Y
PH4g/UGi9GEe2Cmn03Q6IHbP+S1ND4AvrmTg828erUAGUBcnRdFJlGHlxQJQqSY5
B7Mh7kSlMl9A3VhxuKLqLLx0CvyP/BogZ5Rcq0hl6wQ4de9pq9ZhA8rgKVSvYx6V
nU8cl/kZjkbkhHZ3LBqxyUmQs/TVCCILP3dRcGJh+Rs9EAGRzVgFQR+PC0WwhUw7
bGoNzhNQwzOCP5wo3fXgs3QN6Inb5aeeefyVhKJpGT8Beun/aZTQV4CI8g+fo+6i
zEO5tY8i3zVv0Vl6tyM+9hrnvjQw+/AlfPbPu6mSFKGrdwEqfEIyEDA7bt4Vc0XT
BoDhnIAifaIYUJv4LHdLQDd4RbfkGXOWmGQyAASjnAF7QhRQPZNI5WX0PYehr1fz
ewx6Mle0E69wAb2XijYseMDLjWjgmplxNXPY5YBpV7O5MUerRPkNSYOM2EKJWGDo
uWt9zl+sia09dM34uPlegsFP+9O/b2yL1oYM7hFCpqPM0B8PRQkBMLDyclbeT8SD
1W14TEkkHc0XrMKuF8ACspcrfy8NFsTRS1yM0MIFmcKkpcTcDJUxZ78PW70hvNKN
msCppKcNrL8CgzvKUlyjRpSVQ7LTA8FaFkdJkdWExpiNAGxeA2j2nVHugr561W1T
i4veWgis8orFKXdxq4wcOmEg8BUF1Op1C7u8E8MdDULgGucuSnOO/BoArGpVMoo5
PxoIyVfoSW0n/GtDQfLhX3kd/ednVBD+a3xqZA6SgUDuie1x3LInRe4wrtrUB4jC
j8yb6uCURADnimjSBSExdN1S0+1emFiIseMTYbb3/9MgULuE/v4nzTn7e60wYv0a
pi64HdycUjvozKhjlZihlAQRvJL3YJ+NKXW2QM15Czcf6/6S1LRBiNtawIdcY+Vq
fQaJZVWeQawaGqbb1ZRVwU0rVWNIxB7BJ8FEwvrdP8m2XEJ3YdjaJMmE2ddelToE
nrmhIwSG8gd1HY3soLBz5j31SRtNDRlstRRyQfvj4iET9kwgUG8PiG0Qn7OXSJTC
COutqDI2DaQLK6bmtqQubsNfE8IaE3N9lEaaD06IL7FoqkZhRlLTje1YTqwvAwBG
RXyYSAZ7Ul2trw92b1zMgZ7VXCLB3yHDIEkDA8DlIOlOEGTgT1zUV+tDPdpL0+Rv
ZsGK8F8LDea2dYEiiAdvPt663z+sa+B0rFIaVN6lh6Wmjoo6xI+YmITVyQNsCQoP
kuEmFi5BRgLP4RnMusrQbndolq4IPKHu7OSRZY3hoY887yUs0MRJyf5iVfIQ3ta0
4NS8m4VKqEzcGZGx6I/RNCMWuiT2jgpYBNR2gdts2OxfdG9SAiKEpIn0aQsv65GU
vdjLIHQE6fj7jZzWo61Cb4R1qxOM++F99CsRE2ey4Ewcim5aqyPA05QVMjy/HXFm
tDTtMTWi4hjgvtSNuQGu6QzqTTjjx5pm8sTW2N/BvAYHVrueVXowIu/P9FLbtG0X
NSFYChS8nrENLBFXQZVZ9zGCddPlnylkTRiFj2iU+vIeiNavkBZfZccZQQlwD/3f
of5cGWFpMDgh1FEYcjqPQQe/gnrfp7pwBaE+4nPQVR69oTIfAZRREx6tLMxDQAem
iPkIRpv6+PORD74lR+4VQE9lqBJy/eGQrsBN2VZl9dnawhpNmca7aQ5FkCkseJw1
s3Cu2SPwUhffNiJv01zBI0bLvv58wUH5A7RdBwccXZ9TcC+3/PY3emkJH9JJZlBi
eJ5SHvs3Co9862hcJ1nea/amJpvWUyrO0iB810gBHV3o273crsImJO7HvEwblfes
cxhdy2vH1p7TsLjj1LPYp1/HemQr51u221BGRwAmtDxvXtvrgFMh+avKMRm+E3yG
OHh7JYj7JAQW5DLIIXjCeluKOaKg8OVpTeDSljXHx9hDAKbdGk4IZ2i+SJ21+ExS
WicmmZ5xQ9ayR1nJemHT22BYNLOQMab5zGp9Qt+uZxwr3JsGyvvfVv9QWXNFSVrT
Os4x1VPsYVA5miOXBIbGYTLicvOFxMWGkKrQ1pvN7F4fZhsvqEi0TyHzIipFmwUE
F5rQh0D61TlfSHD9+a4eAj2T4xsjVOeTIwENdgnEVsi3oY6u5ahQFDWdYht6bFkd
OmuGXtJeFM6VhAvyWW/K6saibOxtKzcQN+B6EhY7rhug4Nntw6sihCvfq3+rp/t5
kcZcMNC9rCxgZAwtoHCiqJJCcv2ayYQ1VQaIj2f3xVWe+wCAM0B9noxAz7367Cdo
ORhP4o90RKctt8WQWe8mdfEeNzBhNsTkYoO0ZJzeaPAOJXFDvOBpkpW/g+30+pVb
n9q+o/kXTDwPDhSe8CkZ0+4DilBpbGzmdO3/yXiaAMNNC5RyrfzoPoqCARRTCSga
4IqOn+fXXfiiN0QMFtXyZT/nbKWfQpCXV4on5H3pMLaOtqJ//8UmDakekEfG1aM1
wmzsfCe/D7vC7zdsy8lN+C9YxeNyuS37uweEYaz6HaYyWktV6MhKYSpEmkV0QgGZ
Y+s3RbVsUroHdFOorg/Xi4ljxJEUW3eaYKFenQw8nVmD0XfppE6nBqvbkhV4xu+v
WSKVgxxEQZu1iGnZPwmEMc1Z0y4mbHsr++CoyuBL3McpuCtVylfpG1kJLrBp4dBC
Indev7xny1nogn02/yhluDlWSk4zCR6vfufJNs4uWvj1cl5ORr1qpA1zzs5dqN79
fxX0eroHBIT+TcogD34NHzvhsD/zI0Us2LXQJiZVSLg2eSs5DNzfMILUF+Ouw7hc
R/wQXj/3D+6uMoeAEDj2NtKICGKm3llULUdWfaImcRm8ezheaw9VofA0MzYaNZQb
jGdXmJ1icZbm1iPHNRNx5gfXR2sjozD/TrACdp8qYIT9NrqJpbksXPqw3X5orsdM
2A9U/EtNySOwMoWUflD1TKKXPqJda7cFOOh7slTE7jJtn3yk/4QWKt/iQcw5Kqji
s7fGwXK/fua5oLym1XrSaif3BXnZsXU/p69xNUAhrBxnauWGjQpBw0A64BDjBJki
fSbDUAteNWZDHBzVWFtr5qmsL2iecG6v66PRYdwaQJDX5Rma+3HBcBqw//Ymkesf
gxljDM532RZh7dfaDRZkxqHCz0Bt8XzWyD6k92+Hfd+4cSfeDBLeXKc5XWN4dDXr
4HyEuSXMUkRkw7wEZyOV9GonPXFC9LFdFM5ywKIzTmw6bnzXxiwvILo9GwkWRK5v
jmP5dkjW+IJ3k4UMODyhY9yFkkpSA0hKSeoQR4DRBJLV3CanCncqkAMK2rEC+uwd
uzr0xsgUTGWUw69Tc2kjRazagK7g78uGGfJNupCyty9PHBp9oDcYxa6vVhyB0z+N
ikGo7ppZr0wk3LfP2gGN0uwEdGcaMBIWyFxMuYWjF7qMKHPDd5s/TpRNgsdqA6jk
9BdC9uzcbwNE5oqP9Qxao+cpMU/LT8BIY2oARKut+hG2X95Zh427l1lSgbqgU457
3DyCyfCb3s1OxXsg5piaQIjMt4GEmxz6JVi55t6S+qSCAMtRGGzQuYNawJuDu/XM
nRiqmul8qlXHwivwiZkFd25DERMfh7uZPdYMe1xtbPnTvOuKH5VpWxaVFhJMQ4CO
QmEiKKoj9w4lf93xtjn+/a580kQZ9PzCmWW+XjZsXvNLP63Lyu/wREJ6T6TWGjt+
FZJ91w7fSiSlObWD5migfgQTerE/1Q4cT5OA7qXhBd2AHdR1RjnKtBPwiraSqXBn
ZpucyLC4bOGwFwouVBVlfjPMeb839Y80+BmtrdODSzaxOj8DfwT7SbhQ3tIHGtaH
psLqjWEK8dui655qecF2atoRpbl7wHA2N59fwGxBK5U5Mc2RRXsvX71GO9tcr27W
Od8bIngXd/GMMlex/i0mr3NFxsRQhW79iuafGOIxrk1iEytC3RmWy2mAGgeyIxHU
c7ZTyW/9y4JWABgRaHkIfM1NwKelIwtN5U5GokxbHAutKapgqzQvlm/R+k6WdiFZ
/q3CJvAR6qJJ6REN+ELBFMtH7oN6pxctY2/I7t4YI8gxvQzPtlFGoT9CXmb4i6/X
a/L6wAPzaYvv5o7T4vzpFOUaQbfAQlxBw+i/lO+L4MT0/k4rL/bWY2l7jQN3Sczr
njIf0W2jkhwz1erdI3zUPdveAsEs+6N4dywwnbpbIYV6QT2OAUB2mqIZnYXmKa6A
HFm1lD/3v3HQIJYHhWMXhf/GO/wR0cyasZiUHmB+LDpIuRJVDp/73G1uwod6s7vQ
pAg8h2HoJZwW0snVNXCoWAnIlwattbsstMvCd0qYMCi8FjTWw/WH+cZ0B9vpWdL6
i3JwIApzZt6bXt9hwkKrNOinVZv78LUND6+l1l+PaIfi6ywQsFkBNJuF/dAqKBkR
ka8ab4yVcGjyHmtFjByoIMMCk8fixMIVZARWkPYuKvbE8KNqjRisTK7bkigCTNh8
S3cj19IVwX+S60WtEkfS7CalnrJTXeEUrceEnoQWxRC8dgW/oabYpnLsV5dsOWK6
2lxsYo3UolZmAYrGJpOXr2VOoixdr2j35QYyJ7anAW7HgYLtxGUjvUq1AJ4WjT/b
HUEZWB2J9nVcwBbfVHv14eza/aL3XQVuz1tcuzXPHGMN0R9z+Ly2MRvSuAOdhBRF
KACBePdcNFac1ssASUdfGd81fjxmhtpBaMx+GPSFpJuDytHbF+NV0zbYUq0oE2WL
CX/QxedwPM0Kf6rF2eW5vdG50wSpRRXxhTiWc0BU1mDFuwcv4mxOjwmPI/929yXG
+Cyj928pEkUWmk/8x1zRe1nVV6pOFXh5Xj3BVl/611X+5UiFghgSdm3JdehpOjLM
7qe/q7Yc7t8tU8tDvt4tfvDmL3nAlhshlXyCe8EV8noEFBMxHbh2IDAQIP8dzUPl
8TfUsNDHy/8l0kHaPMefay0iBTX6BCas0fFDQvAa9vN8JJyfG03Qxd1whTCbSoYQ
go1SQeOtHi7CSOEhmAufETd4i1JZAO3Y+s4CAIjEs8d395dYtKGzsZBEEQo5Yzq9
fWz/tsWq2xoHKZHmcAgZ4ockuzy6bXWf3QYFQNF8tc5kNK9b96H91lfFmlRiMhne
/TvYSHBZrwktGvsjELuNlJZY7wMK17YHvsOSgv+gsdyHmsvnqwrdNIKiL4USUhPg
YVdE8TUs0o42cBki/1LGkQVMZSAKFzZjUNxG62rv0K9Vn6kyNbbg7CTwEjFIL1fT
pWarxZMnAOmUGaF8WPCFFrO/RBeOl0QM8rdiWj6QHJE7WFXfJR3/z1IEi8ySnx+R
qXPMb2p7QaETj+u16ve+GvOnYlipoO5FyT+KUTwfQToQ5VspApAhtGSsbiYg+5H1
yqPFHpqm/oa0JQaLVmgC2PnbArcHEFSMxJdlrSd23Uty6TVf7qRQvvnwKZ//Vt5v
C/g4778SgqFSSnO902EvhZ2wxZgSJY/ZpK6wMcTSc8ManSXif3toIdmHIbLXbcSR
3xfSi3u7DpeEYDUNI9npHmCAye3h3BFrpc03B6Al21wMxR6A2r2832jDhzrbIIRh
gg84Fi3BKC3GCZOw1x3X65U5oRzNqlIKp5fPDkDHTrGhf2AmYZJFxjRKQtKWY/wA
NFWBKkQ9ICgG7Z0oeL0eFmxS8kkNHYqNO1HbuhMalm5jVlx29/c5ZAVVPLci//QO
JAHTWGJulcGZh+XXEkXwzG6XhONDrK+mMgWYKPCLrVGMn7WlcU9lDW6rPMzn6pLS
L3d3OTJq6b2PnYWIWUUYTlGMJDIdsnPgn3tAziMPR6ucv5A5NYrt6lli8WJw4xp+
D77zxXQAhav+ZVbTtkND/Ph+/NNul52a1LJaY2bseSQAJi0vSasrvm/erQslb2/E
YL3gFErb2HwbaT4l4dDKBnOOlhR+L//3CxZUy3EAzh9XUvflpepMA3XkpBz7eQlZ
o66Wu8JQgAz16iOS+h8gBRS8vWMx73OoP9uYhN/fSBEtmvQV2l//k0ZejJI8cGsZ
11aFvSAMFFyzxbkXoP8Amr5EnJxofKa8n/vW0vnx4QuCSzIXJCmD2VI1wELIwHL/
dgWKpTo2bOaNPl4YvArX/lH/ZoCpcMRxUqI+4GnihO4Zwcj7mJGAJJ8Ng+wecpz9
/1EBMO6bnj5wSmmfvczYfvBmh9ohROWKWYo4ebluAcuHunqDJPvLptEahZGZaVrP
RTdz0DNgdl8tyTW25wLzus2HABnDjfP6BEKLIyl5KhbSLAO7AHEAQ2A1RlZSwib3
WWxHXd2uuSNTSg9HjMWVc7BRWaGVXaN0lO82rsWZPUE/TlqCxSaJbDAegl7yGgp2
rsRdxwpIL1rbo0zSSxv1T2LoSqjvZvui7PbVxzPZSigc56D/RDTrMQFcaFMCwD50
9BscKJ4labxKNfRN1D3LHRcVWFr1vurM1u3D5z1UgwavproeK/CT7hXIYVl3vUw3
GvNKWu7cMmSeBH8GvN7IA7Utlzl8eGFJW8c/imWZ9kghXuX3BlRkSwtInW1hophE
JMVdvVaaG8HbFt+dIZ4zRsgPRgO54DpgWDkJgDVZAFc4t9Ls0Sm93hO+YFiJWYNE
S9MvSPDtXQqgck6mefMeXIKGqieV89AFemu2fsQFsaRg0+pezK5DlBCiLOrQCN4o
Z9zE8Gv3bh2etRxXl3qrrA78nb00x2jUUxFjc3sSTkzKKQM9/NfeXGFXc7QMFBdg
mYMlZVJglEhJGB5xxXOG1xWxjbgz+m1iLctw7JpOAdq/hrmEETNEEbymCvOf4F01
lNwGkW41GWYCVdwE77OcprlPyzKIWRI/gUJgwFSiQ8mQDCirJBwpvDg0wPjIjQts
UnKC2gbn5UCZEA/qq5OW59FoPdJGzrWbyXgvW91pRF55Q0bD3rYJ9MQVVZO/gpnJ
Fk7mClklLeZkwjczoHot0iAmIjUpSj3Q12qaArfxC5gbP69nd5LlKxBC3jEXwZ92
zGXnBDGaqJHeKoXRFVGrn6PZo57MxjeNAhLjZKUaqca2kkvcKzbTLcDr6Yv/6EXS
hhM1kRY6ntChsQWmEO+iyFAoxLGK7MqMXhBSeah2tiIDqo7xa5TsbcR7xFBnBa+3
rjKfk5pz5Q4zWkcYKl06XOE0fUYHFtmU4+ipyHrh+T3qLf9WJKvtqvZ6FeJWYNN4
9TkV002pbT28CZFfclxN5ROU/q5QuxP/42Z/b4lUTI0xIca/xYB/iivYvVY4LEHE
CCH4ANj8Ix9Nfe+xKFpy8CgI9KwRSHc58jGKhzF0qqCaAi27dQaqrQD9RYpWm4qh
xHtfHy3I7v5sGwnjLXntcvfGpnm31gqg2e/SMETD1okqfSXl/Y6l26PCVgP2DvT+
ds5FTLiAnPmj2D2orLaKzQ8/MPY20eY+0ltQujD47qzlzNnUhBdaxuEJXywTC9jO
8tjqOF29eIPxNRoY84dgM2pRDQ3JmrvmYLy7SxUPuyKipXCIKiL2TtxwMzqDY98P
DvKuRY6+D4r+xlCOktPz15cjQzXOVu6nDZNjo8p0qzAee1Rh/gqRVNgna5zzVVyw
3AUJD8sBn9EUNiebZ2+RGARQQIngr1S9uQWEVNKP/U/SRAlKkjX++r/rEWmlDAdR
ni+N5uSogaq+SGp7CilqYEDyLOwY+XlI3tbwbpuEwgqZFbiMun/Mdgq+CiGRk7MC
pRDcz3uKWObjHwiiTdbk0v1B8nxFpZ1ZfGiUP+ab4KR/nKEcDcw3q4+lG+TRKzDq
PXW2WNmQtC3Og0BPepVXpN2BD9K1D63e+R0a0ktNwOq6Z5YEs2EoAE8dXc6oGSYA
N9d8AbrtGyU/6fkRt/0mDKqW5Aso24SDVr7eJGntSGFMQoeZq/Th4LiZARtRJm2v
HWYkVbv577rs5l0tehDqB2R6R2IdFSrJLq7FjhMs/WmUDb92j/6dosLUNQi4JDlo
QTofSy0FXeCPRMHvDTPsBEgZrYelGZZcnF3C95Ny5d3Fs+73VM0HBiflfX9yugmm
PGhLyetELJ5Y4Zm71JX5TV3BMc5VukGwOr2+RgK7ah5kQ9+3kEkyQLmErVyptoBx
16JruougDo5QBkk1iUeTu2oZW48AkdXfOdPcwzRpExdUiLDcQs+/Cie1+pOj14zo
wSmOzP1PG4kFYqHsDUehLNOr5a7QE2CY6Em5Oov840VFfJzzQ/ogLnoHEsOxf5Sm
KjFx+NjDjF1+tECiBr0Q2CRUD6TR4gFzvWNcwAIP37tl5TSH2Wn+ePVsenqDpNEX
77IG3+cQeXWN/twiIfJT2dW6JGB/UGvP2ApYsyvCZBDkv7VEMfakgHGpt6Y7Z7gu
BolevVrwl5eHfGHHRXUlAPJrcMqstTvG+u41LOUCnigfXUEUPsagpICjdBjI62cl
5I3hbRsNmCTmJ+7Pw6Zccf1xkhg+yNCJr9SE2/y1/7cFBeZyMsunh0tBJBj7CVN5
NFf/MbhoakJOhOdjkueXlZUiw+0oTmBFArGoNmvO+0RCMzhYgaGarKBAaa4jscyC
2IrrfsASCSFhBDO+6KycCpwl8VayH36vJYqfW/ZwT9/I9inWnwb9C40is5qhyRd/
263GvDlvNUtr6nVBHzweuaL4zbS6a3rAvKtdnHxqaDByrMIRjmG82uSn/FyHK4C6
eBxag2t5Mq2XFUsf7cuTRiBeX4jt7SPexZgBlhkoODSvxtYRbdwKWS8h0iegku4b
maz9Fw9KjahwRcRN0JxCDjz0h5sFZxUG/9naF++U+0YKxksFFWZlhvqJJrKdGyMP
LmF20qPjHVeMqLy7BErRTWZicfTLzJFlBzK52OA52YHSl6A51NEjU97n/2Y1bvn/
hmjHHtlhYKFzmoIum5I+RZBjbozmSkrUu7Zfg22CG54VPBobzk4oc0/6QCLO84Aa
X3EPlUfI3t3HGFIXBy5+hgCNrz4PIC23DYvVhtmSQzqyltMJ8aCaDnCRPPrb15yq
8nxx/R1K4ZOWEdPHB6tYUrdqZ77Y1HZo2UCfuBHXp6xFSZGUDmdVkxwuemxD9uz9
Gu/H0Kdu8Q94gRr34QKoiWGrmcY/Up0ijmswrNJujSjd4Oj/CoPSPjykk+/xvT2q
Fzj6qeO7YC+8AM/7PnhBhq/N0v/SwbWoEiceZnJsm4jCCk8aD/SxtLi8/UEw5N5g
+mSSEZNduxgFWFItZ0YojGPWgAF4S9GGl8Lg8S67ebiNxyM9jebZg1c/QfqsCO3q
qtiW2m0QLRQyHDUlpicksJzexpexS9g6vLECzggWU9XmWmWC5Qfll139+0O4Xz5L
HTMr4/MaFahLhTCEmQlg1D9OLYyjvvsC6iZ9TywiV7ZYgFa7CqATAUZt9wvo1sKv
3txUdOs67dU9GJMftQwPLOmwZF3S4uabyqi6685NykzVjydHtvw3I2dEEI5qux9d
+aJtWOdbClRDrLj/zlROmZTxDu3CXJ+9oAXy/uGhLw6qMZpzf6doBdLHSr4vCuqR
Xq1XzG1B0cBWK/YLAGoDL9CXk5573WSL55o29MbLVZKB7Jd/l3sTehJz2XFdv9It
RR5oGDglhpu3FjcChkBjKyz4CtDw58W73r8ZVFwHwHH+KMd3SEbFxUIsFJ1n/rzH
ZnH6iexR4trT5N3vXvT7rRTV254caIWRz6R/exIDibLqvA9NSl41tVXRfZ3L5qMQ
WdcU3iUr5BXQYYbpPG0eAnrLV4VGabELyKYacwEZlZlAP+Qtab0Euyi6L/e4W/D2
B/KD1Yf+EpDykFeZV+CpB8HJldqvWPD9pkANBzDGLsFXJFQJmRSec32jL6Zl/WwH
MUgKGcrU5zweBB/4X9SqtqCMayCZby//P2xyItZhWg5dTNf1+TOgaofXeZekzFb+
Uf9dHaz42R8kLNX7x476XXx050IMvgDdN3RwgFU5ip32oWUlFcbDdM5JYbhJy4te
d2ptgZhy8LDPrjRTBVMDIQ7mRKr7Fg4r9KFfiIDmEGeEmCc8SCm8cEbyLH4M7419
9BHwbsFY3yhOW9roi6auWHKSG1dZfGKGrmf3tdDnQjnolTV0svAteVI5IaEJvtt3
U7+wuD/D/zFPHV6FLNC66YhcadcCUooSHVogSOSDNJ8ZtFhQkXESjdUq/g3bqzIW
sL9KejqimKWe3YfQ0NbGQVgSEedrohm81MhMiCdneNq06l+iYC+Hfg3JJG5lOZff
x9u+2+lRfsmguX4WomJxxn36AmKEhlveeZg/r+0FoTLkWxqCxFf24zZNTH52ivO/
39plTNycvSfAKX1y/7Duos3mm50JuoMCt7qydg1RqfNm1Ws4CwRBLCzC0R02b9PQ
V0NoydRm7VuE8SpoZw2+tIPpbuVS95S0So3hNPjKLU+Nh5rSLTn8QOjsEk7pOhdY
t7FDWrhsFupJv4CFU9n2xNmMzCy8dOwrQ3YBns5JFv96noPdiDgMouCD7Xb2eche
QOxujSMqs+yQnN9hPRLM+HzcF10q9jAhZyC8XfV1i3PwF+ukRRYkgEOA6y4M3bZs
sEYGRelggHItCtEBeKoTRBI6gU5b8Ub8WXTGw78fsQeVgAL8ANArVB4bNW7xK6q8
RSqhXGrSOZTGOLVch85sKuxS2fI4hsILcSAnjuK3Y/VnoB4/SDzAVYnI/myLxEHC
hrE0bwN1z6O70soEFeDL2TRO/woiOl7MpwXcyVkLGd2lUtOMA9f2j1dWjTZr+Sgn
pawiI0+pmLHnBX1mQlLf7JmzCwCC28roY4d2x/E7ng2c7A9tXz+Cv+nB7doqipuK
yxuAVGnsxOydvB8bGREAvlJZYl3qwcerP9dptMAe4xxN/1oh0D3zIz0z1x8sGwUh
H9Q6L2/9mETd0QQ69/PlWdfFuEVGZ3h5O8hJV9z2Y1vm9cOrKmmB5265UjImzt42
1RLamQOy8sLDDW6jKraiQlupdf2TIkMG9ZMHazv3C2banBHr5khEN117/iCtfwMR
wbwjQ7RtBy4PMft4ekTMM6ZMmspdeQMtpcOcWPSG5P3qLirlARk9CvBD5b2jIEY6
7JtvRJ8tsAElEqRNEzY/ZuBWa3PMqTmkAedcsqTbqD9Rcwi6S4q1mhJtg8MRT+HP
1NsLtYvFplEQ0KNqB3DYbxbojrNyIacVAu3A8nnu1QlqMCTTfk5wD+udvs0nJg5G
kN/bFPjMrmxbFl80aTFsVUPYG53jlZF6PJvA33VOOvQ1VfnkJkub+RtMz7ABNmEk
BJtnT1SI5E1QigvYYyxooIqshLi6bqTfliHLKVDooLQGvWwXEs2whOYtYG7slezl
t/Hxiq980QsI2XUa3MGpMPt0En2QBXD2vRVKXBxoRxEmJTOrDj25UjqSDGJaXk3N
EakGOk86uczRlJcpVZP5eaGch6PsghR9zxSz78C9wGqpOB1owNq2MooaEtsmZOt7
chYQgkm7qUqkB25rSiJ6bSUze52i+pFN4PpoeZrCVZbHDLMHU69mGcrOZScYmeQ/
ZlWhGcwjmiFp+QAeTnnX58erZL7ywwProA6dhIpEPa4olE4iSZ4EjH36bwnYDeMO
KlnVBvQjkJznAQqzYGs7eIGkK5+HtigxPpidTA0tpeQ0jTXoqmhWNOplhdp+zvCY
7oe0bWlQOYPjqR7pIwxuZN3RuG9uSwMRuEHq/P81MUZPydOPAj1CDDz+Q9ge+TXb
jzCy0jQjv3D7LUpDceIJdTNXd/F3YEN4Z6F//UMHiZBaJ96LymSoAXlrnTjxlybh
gkfDjapA88pWVdo1M8XzWC76GnA7pJrCL3YSK1Wa3p3AkCL+wBfnqzT1UT0/dJ0d
YvWFGifw+L3MG9n+3KvL6WFZuGWKDIp9VMMXjYh3tqUceDkteZlHQyvX20DkZQ3t
BAdKZNaECL0TIM9Q9/5Efe9dnWqZk3sCXiMkz0ooEREJgsPfw9p9LNGB8JVc69QS
GjHQeYNFdWBlOeJy29sTo3Oj2Nzwn3T71dMudvlf5M3o1aUDhU0CRszrJtoKXTER
dMAzV7SpcfZpLw8bvupmQh5eCzT/KYMTNunZ2/dMLQkl1KNy2YwRoLEQOF/5SNhb
gD98dtYns/eplvLSUDBygUBk3fUsaz8AFT5BlLg32WrgshmrcQITm+0JISTbl/Wq
tNJpYfwstaCBpk8Cfox6ZRIR8oI8Iob4s6436dyVrvHbQlQpD3Hh1TiJyUm2ejYc
osA7iqf6H/VhL5tCIohcnMVgIAjmZ/qgsipT0A4Nd0ntOm1oUo07GjSnNhGlcESy
lQcV+02powx4TXE8xt/Fhxgk7ibZ1VginlhgLl/EZAFtIZYzflMaJoLNZyN+yfa0
OBso2AmBMyMZt2EY19Zfduc9EHI+GMaZOzB6jx0kb8qpZ2ZIwsoEkY79KpXwZ4Rv
P3QWJ1SZKU6GlO/BQqOkoaWLVUGly5U5y5Q8yObMzdCjShes70ZHlBSDg0Kvijz8
NpyzruvpIRnPoHCjCBREzNu2oZY7g4dFs/6E5ESZi8RES9d2avSujb3CHgNfhu5K
/KgUFC0fPlJCB5z+evovWoZYhNTf9EuC4NNLhmAqj4Totx5sWao4tYhb9Qvl8fEa
4maWLvf3bKFw/vYQIua2dkf7EIIu6lfSAe2b65GOd7rhkOanXs/jabGPlbfrXfI5
3KpdsHbaGtA0Ds4rhuYdVEnaXX0DGFPleS8BUK742tFtAqV8eklvY9aQB15xiaTq
us2lJ9TGMVNQE1cA6KYwTRR8kq3R2efztKWizRRFSIekPKbIHLE4Nr84QKkjYCaG
ph8GlHyMB0mVm5w1pxKtM4lkMC8ti04RKJe+VjzDfXURLfdFVKEUkGuYzW5XswQq
FdqF+LvBl/wv0QPK8gjpRenpUEXYxnVakV7L5+V7bMrtPSIr4YGAjDGxacLjc8UI
Vm6hlyeWUqXe0k8PK9tO67pqk/tylez/RZm/6ux4sjbyGftdZOOWTb9x5HVyS/PS
BwE9i30tJdjbEte+GLlulrMcHTDYN0jYjTEe03exQ952CCXYNemF8vaqs4dMrzlM
oULCb/LiUy0wY5lUD6JWRo2biuHtIuotvft17ATJkqXnpoq50IYz+h/RVE5wfTNn
sJi3u9Lu4lXXFdiaFcgvP68R5tN+T9ZZEOi+xmqmu3FXLFXj0d1L6hBeRsSay3uw
uBJhE2n5G0u8pksBMILe81spACWVaE52ZO87Xewa6VC3OqIM4KHuYhuvfsurzNT7
La1cSm+wKewWWU9jUfnoe+YUSMsuBnHQYVUad6apzi/QzLHbL/ZvusQS/yVWetn7
Gq0jeGxyaZV+cgAk01BX8uMNXNDfE1xhT2EbQ5wwMJWTkzcldVVqTZJOqZ3xfgAs
AXP+Chu+09EalyLMs8ncUE0kvvGn5d+s74Z6w7wZSVDvHKbEq4D45GAMJnUpikvd
vRK3Xffq3M7t4JRzX7gBnH494zhDq61Phyv9biBCQ8Gp/l7F3giuzqfvA+4wRD2q
Wgy3C73SoxoLE116/42OIHB/Ab/ZUE8NL9/JXQX59N2rdFcEFv2JmLKjQPuhlDbh
StOpsqtfdT4j7jVLOS2npA6YZdWHGPTDk12A4o4ly5wmbqYbIt51YsrlFxvy+qpR
+STaoYj6SVWkPnHKEA8bxHUcuIVQUFQwi6jML4DxmtF7wjQdXhxm1PzhO4JtQg8w
kmT914diSlnLE1XvnPU75mnh2kky8Kz1L7QsNxpIkiAQHZgGE0PzYcPq3CLu/U5e
EtldM2grc2RplXWexWH6iD6onCIfojsBq5a5HRFAAHQ7HSb4Rn75vRMCoudauJkS
ahvEOrFgzQo0mzUljtPlUPpifk9r7YJZ2naMoC92cz75A0L1MA2e6mHIFfXSaE/6
HCYkkO7WvyWO4LDxJFgCVRUVSZDEPm+R6JzI+DfCRRGZ3OJ19Xi9JBgBfJvrgwpm
kvctoc61HFhcG32Gj1CzpKEu2InFwMK4G0cuRZ+DFDPlT0IT+5H96yi66ogeFmBR
uBPtNq/0ksbBm4RJsrFLaBDVRjrRmp2JMxLt70ueJ6EaFzbRQRzZHO/9X9XQ48XY
r8m87zxkuH/G39WFQgrXxnzlaC8ZNGWyN9cMq75QheUIPfx5nMJtbKdBM6qyEYsO
CCJH7myXRIj0SZ+CKZpO5co2BkybWW+Fb8ujY1xwJQXVBLRpr/mp+20qDuJP4j9O
Y21BWqZC6pjwoUpzqoHg2lDkAjvmHNAvnnWR2SwPDrDkTnSMBiWa4KAQimdHEYrf
410v5DWky2SxgEtwKSdYee1y2L0IsSR6pPvuXs2WV2dZNKgYf8gpbHZIsg9RdXB4
oF+fVFABRio0ye8eMNXfMSZH5jxNuIxABX/b/8JTdT5WoUtbTz/uX8NSPeIlLLEZ
Tj050Repz3IsHyDh2uiDe81tTzg3WI4mjTRNqjQ1o0Wh9gH3DY5/rFSjDBSOPzTD
BTcuxiXICZnSaq+aaVbdxySnmUN0N2RRvqWYbpnMYugA2MNqorV1pomJs6IDhws8
pkNmcy1gmCRw+o+kw4JSgtf+aB5xO+ky/SBbhgcRhRNo6fyAq0PXoGPRTeYtMj5q
Jb7j+5EzbZjuCILmi7I8NGCCswnij2hbcyZbu3tQ1QiSqzqjwwiQHCQ2lzytZwHd
Gngy6V33RJCT+izbC14tF3Ev6Mzi5zQQKb7MkEKOQzBREA529uTuw9z8qdoVyme1
4tOlN6V8vhf7NEo4BBY4+mSSwlvoHd1C7cTNdVfLIkaY3/FXH09BY24WhuxTr+D4
AYiK9+volXYmoiT7ClwDXJ5+GyTQNH9vb5EOkN1Lqd951ByeStVYAxG5JPtM2AOW
TzmoELhN4PI/P5R/mnvFkewmXM5191JEtafH1qd0FszdflrZ1HQdbqkutjM0f9L5
OqxkdZMFW8k6XH25oyp/LmOtWIqR1d9ulj6j3/EPtjOSLX911eKRCUZ6SX01ATvy
8sNShLhrsJGLAttozXUWZWMyywtIbtXT7j9IPt3dZpJEsacKJVVTGbxyVzBGd9o/
wkU5SyHtNWFDqfJJVXX7W5nNgXyodVLh/qFQMhaZuIjvW3g0yaTQz15/7QdIvsLi
XL0N2avoNbRlO/9ZkU5iR94ojy1796s4xmu9EC2H8GFIjjcn2Ge/f4oJ9yWZydnO
TWgfjnJK7An6PiKt0sYknY6sHDIzMHIuc1To7WThzDFCsOb7XSo7DhtAjpch0ade
p3zjvtqOTPE3BDwKsoxFm+abRocAaigz9+aETPhxDa94IUFcoYSxL2VkdHtrtV1K
5og7Suy83lnMpd6B0ptmRdwZpx526K1RFbCUHrB0n/3Fd3z7Ed7dJDHAoYXvdT1T
gjbBpu0OlXcyAzcxRDE3AgPNb1eGnyJ/uqMQ2vcMO7HQZdLcWtCSXsLFU5nqxPsw
srE564erjLK0SYHCJP6vQ8d2F/a9Er1suhD1TRSvUy5pcA37MV/SQ8JfYpc03h1z
A1fjYbZw2WPZSTSkQYhbISGJTxKw7QEyZikVISA8ykA9mKfbJY5e21cb5gV9sKl7
MOHwPgUU8pm8XjqiB8OGJ92e96yZFR8R2ikDzjSrKImSBBDVM0oCiinMsS2+8ROu
c/wJ8ULT9gHwXsf+olKa8ZVgSNPPasH+y/yUXcBPQKjmf61s+CDD68syPox2AYfJ
dx77sQ1TwP0raPoT5n0BkMc1cDqpqvzxicxBpUfgduKAO38eGD6x8eOFsDzzBW5g
Qyiocxn9LNjTa7r8A8wTIBEjz9LHtfEfvYlMMricbAjKiHPX7SgeHqyEPh+Gw8bf
S5fh88BXkBHghijNJ9wgIOjwZ4rNDWIgaePjroXtwbS0WUnxPbRiCJY3JY3lFE4Q
o4dTh6wy8WDE75pyzwkjHTm2h7kZZqzFVAEZngZNxlLXfboz0ik8u7dJXyv/Ym9j
x49Ql2P4p3eKMc9dGQbutC4yQnDsEmfC1L0vcyZSnpxVcYf0Xx+wevxy/bhejNKE
+x0La8S/1gqrxwCIWoR8pzb8PGe6LuvVKMXPlkH5HbLhA+EIQP2IwoPvwv19EPuX
eBlBmYby10Hc/TuGkzdE/USCg318EjiwwSrYHbUjHVELqGoYtX8BZaDKYXtaRPN1
UTW+L45ptu9BR3CQM9kCYcYP6SWBXFA755xbqQeQMnxnvtOq2//gsVXT8qU+rVz5
0IV4/8JmXy7xMvOvhLuW38ykkJ48Cdq0Z7zne7ITFh7zn3lqEVJ9zeKaOe/BR97Y
vO9YhbB7bkMrHyzZtTY158FsM6xgdqPeHed3PEvQR5FA0CEw7wxwqhJoguf+w8Km
UMAbSak9D2xU7O0SiFVcBhgCU6w2mjcSDdr3GkCnalGQztjmP4h8pWKL60A5KBt5
p9U0ibwa/5z2N5p4NNRdyP/e9RrD+pz9ist+gd2H1lQf4BvhM6bylM7GPbw8Sc91
EiJUvMdBBawm2a2C2uXH37KccjYeb8i1n4VQCkJklzA3d4RdyEPrnG3HXaem96ae
3HRHFGEndAyey7jExfQIHQY2xCujb9Bxyfdm3AROmp/bywhlOIqbCWzuhDZs8fiz
FWZTzYlmVAKgDjNNn7Epi0gwx2ktWzuobyINBS091/ldDu8IAGEJCaDJMQayfFHp
GXF/ePgsATkSbfCTWPUhwL53VpP1dCWkHtid0RHeVTQt0CrMYkg6A3eyOPI39PPP
I5fcihgKb6y7Tgz5YiuVGZx+GZkxm5F8Mq6IX5Qd+opQVx8tfBhHjbgUeA+n3GVf
F9Psq0JtTgJLEUcDcrOLlI+RSU31Q4Ld4PWDS2+4QiU7+30i6FzM90NJ7+EvjcvB
rq6K6De2sQsCEJrcx+7/5QDHNvyDev4AIxakKuWMQDtWDLu9lnI51/G27D/5aM5X
P7gbyXkA6HxAWdo20x9X7fbnyvlzh2Aw3MsF9KfV5WwRLHfuevhImfes90rgC5sd
vEfrSv9N4Gn5elyHYaGUL9buG5ARFybkShWChaRlnW1T4vQbQv7O8WmcIt8ZMue7
EIpGbh87s6KsYf2QG216Om/Mroj6BIY+hTci5tEyvwGrj7s4m3OaaXDYrWegpVhV
UP5GyGDans4HGdOip+O1ODrd8sjqCVyjDXLNa02tiay2MHneC4Hj8D4k22hhO3Le
cfo83K9ZqpkzQV5s4907ss0sPQhW0xw9iCCWF8/CkWgok9tbtlCPzjPGjyR2wiRR
vU98prdpxDusTqYRcEJ0o5cXlhHo9Hj8FW1Hs54NwgwJKRPUyZpD14QNK5nZM8nV
yX/1ZF0RP+IeBAHLh+l/+r7vKXI7418AQCfROGYqjMzjQm4Hf2vXKSsswoUSQ5qW
fyXcGhwSiRT5dNzLboUN2g6u3K74lNU+towyFfxKitQgTROx5wpvVQ6fxDW7qVJD
UKB/u5vCa6hqbPrq3TCiy1IqkIxt7FOKFg3cE5Ad5lm9p1X9cggU26Q4vsyUgQ/Z
aSU/2GfJxsG6br9q1azqvjFM50Qeon93Wf4QWITPJVJ5Wi73rHP6F//Xd4hN3+D1
LLZ7V4y9VXkXwqshvAs/K6BsJPeNikGbce4Jw48ByzxGZjZrsCqVkFuDIfAhhZMr
Fr8zf+0fnDVk9HAOY8BIMZDE1tPH80hxVVyFOjNp4mt+zky7dRcuYLT61TcA85wq
njID2OWCVd9Bau/7qZDYIWf4IGSDTH7yYabNXYHDMUfzTeKwhiddTyzCt+sf1mzI
CwLs/NALzjizp/mzIxrmQdZuE/OsPy0KmMTxf7hkzv4bazj+4xvdgVgi40P87aPT
2bkxe5KeYcQAABlrgWD0/mYf/gZ1fwZTd/4ZhGa75YZv4IeYdBvHI54qeBk6CUZu
E8NtPSm1P+DJJtjVXx5d0jZsH4tPPnRMVHTO8WIHsETeSHJTdaUo1aGsHNiKuBQX
avTrA1+YTkzt29jIh9unZqF9CRMb58qpFIMUlVY3trE2jv2UJfR8xj6H0buXqJd2
uzFW/oYIMMi81dVALhj+7Lh9HNbTVhozI9/JXB6hX69lbOIWJZlFtJDcFPEHziuX
w8+ncdwiqqnV8AAuROxpE64MFHG0cMXQdC1SpsR+AspBxj63jZuxfGd6M86xcIvY
n8WyRZCEwn9mUAB33slT9J1WYzavCfKKOzTeVmUR/4/fLL1mV9zoLL2k0Yk67pKk
2v/zAzuaEINT5z3URZUlqUXvKSORjkX1pBqna1VS2m5iwAIoBWZxPQALT9C1eiPr
fdtWfQU6GpAlnV/d3kR8aHoel+6mjkYwQrG2ggB8Yyu3yt0mlfKqEC0H876Sop0M
3vi7at4X2Fd599XLYHDQvsCrk4ExJDORiEDPpx5PdisGobxTmQDP5ClozaRIdXZJ
DFaNP1HKApsS5rpyxHGauPenkHYqy3bX8g8RXtMCsHIL+YW3pH3gogDOeTT4f3BT
sXRfq60yDG7P4p7Hzqm4lqLptGX1MCYcVDnx3KtJ5snZn6/8efJT4QuU5o+KkFW/
SYlbTl/+I1667chr50BuObvCj5ampEnerFEVerE5EnETi8q0OY1uPlXF7WmvlOlM
e3j0l8Dfkw2oVzNo1HTe6Qn2/edtk67FRi7TyHKCONzS2fbgwDq7DS2Gk51ygr5q
YMMJvF94OK6U++JfhGLzjDb+kbxSr69OCcOnAItxH2PA7iKa5jjTWzfyo1LBrFA6
dX3zKMRpVrk7sryw5PzRseOR8lkQ0ldxFpU4/rB5vJ+DWPwFkfXiklLbjBkRZhbb
LESbXvPgXEnm02gV1unGMNJG5CflH1oubQ3ol2nXHrmojbUeGo+4+UBW3gCT7/Do
url+EU+/5a1gcEdf5OijZ5ysKZte1DdLyP5i4QyBuluzgZolIeywmPO02FJsxz3I
0Hf6MeO7fMzZsKbHrTgF0a2nH7Mz0NSAbh300Ka4ae233AqKXtCuri+x4ogpV7PZ
RHhvlfWauVK9h2JURFmsV+sykKHUtinr/SIRKBBEcXkTXDtBny90GNr+oNFE0ZWK
HM7yxo0AxFVWCwfj1oq1gW3lPyh8lUrZUOVdyybUO/UDTwnQrox3oAljl7aadgci
bmevGYld8JI5dZX3BTNG4Rz/QcaUhynGPt8ZJVHQoBqFWInraU37T3z0s+f/W2qu
rv21X5w7D/tbiqgx2sObd2gXbCvTKAG/GvD0H/hQrrqqEbfevPws6Uv/+AbrmBiI
fwh3YhAe2qEwA8CUi/wf2pr7jffWHbb++pgUXn1WmZZqC+6bCiJCYeRBU2uxaind
aPvM+3WqjfChzkgVxXrGqjP2LUv8eZ2VwWFsaAXw12feJapd6FBcaXPmfDjvKnq2
qGcYYudVKeF7HCWwbFZvtyhtt/BWPrCTEb329EN9C/MLRykr3c/yTbgkN2ekZnZt
8JUnc1GEjGeM5TjVcFNJXDla5tCBQFDJrmcCT6o3p1XMrJBQCOUS4uGwvMH3dkWM
aLSs8ehPdoAJoGDuPmisc+1ReM8UxlxuV48OdmlVD1iSS9GSrZy/N5ih2mwhsDW8
N0GA09VXhSCxaL0o3NlFY1E6D2IhbB6krQW4U8y1G9nsX1q1DiQYDlvWDKJn8+Dk
LVFH2zUuzGklqWeslgUlzidowVLmAxou9ePnwn9ERSZa1TC3CujlI9/W/Tovi6gr
d31bEXAJ6n/9je3VHE6Po1RGjeXnZJBqzcmnsfPHL5sCyvkrLJsZ2SRnpfDEIhJr
zRIQej3Clf3psAzfWWo8uq/CeHKI5n1/N9Gppc54Ca35C0Po5BT6LzMTq7ZgmNHB
T45yMbC4D2Y1BCQaaySgf7yg5rIxudqmDRrKyLJr0NoyQXNfPqPV/ZeYpW4H4bI3
EYKuBvk8FRmtJlbfZJIUjQ2JhJTCf3zbCTpT0QweLa/PLdsFiYVfQpp8CVIdZL9Y
BTPJAfOxoZfzUwoll3Oju7p4iHGLIoKMqU+tnCKjmIYZ9mjicErPwNgwKmgO32B1
gL898IqiSQcL2Q3CBhwK+4QBtrVXkEuarL2reQFbUANYSSUYoshc5YOLdAC+ArrY
EKMZzTMUTbEFJwcwfcCFAAFt5YVYz5YkEyAXfnyEcF4TmWaTmp9iLMgzgfdm64wT
ND+08eguC9egNrQFX/F3VzEpJn35hJhqB0BPW7ym3OEp/GozZ6lZRd38vi6AvqAo
4c+tlGbEdlpu5scEc+rgFJWdTgGWF3Ak6nsRsJSVE3JGKHhJu7YrvEpF/iLU+iQY
ve89bsq+por5ktGUqeVIBLoexEel/S1cwD30tc1Yim/rZxpl+444XofIh4UxGmmS
JoNQUQUj/fG3RY8RDzOo4Gr9/Z4jlHeLv7A6A4qpFK4TnM7nBeW9Mxu0Sem5T1Gl
cV5F4fSO6rplTBX0t5RZhyO5BssVDH4Q4jEWLJ+6DxCHvNBBnIgVPWGIfRtqt8jB
M7IrA4M0r44DXtlOjVC8Gb9ipTB92HkkSxBoaBRtu4z6/ArjPsgCqJCzvSkkRIjA
0gWGpeFAXd0i4DswvNTPlmFDEsFVLrRlJojKSufi7+1t6ku9SIV9OB0ak5W2rC1o
dEx2qGvY87HcLEayHX0d12bJYt59FMZ4OphjboyWgtpp1N8TxUK2pnkCszzU8GBa
jgyBLa65SffemkpeQ/dbOq0ZWFB4UOe6yo+feqop8IAs6i0eKzLBFjYIdS8qV2Tx
9GB7o7gyInqmE5F8xKAtUK5zXMd+hR/VIFZ8EXNsFIQJUlXDI8A2kbEHhRsoKpF9
qxZqVwIgmRBxZuu4mTCPB1IvelKu1+yH0BPwBlKcdprfuX8NFvhFN41UzN8YeGwx
YP8NhDl/hFcyV7hkpI4wntxbohwW5oBfXflzNgn/BxRp5p1Orr2ePNDYMQnFP8LZ
Lu5p9cYLgXykRDJRD32AaAL9exkVumiW1Ba8VaPoXfK0PxVSRb7Q/3sE1jYRi7qK
RegAgNN5J6uopfsdn64o35M+HGQeMNHIWs3x5S6AZKAvvG3B2YNChae2WblkN5Id
oPguCfRv676EcWCo5e7kOihTgQ5gJnjTpRQHhtGGY5W1ajTtU3WclcKX5TzQVnnl
UP0FM0/zMxH8C9zXJNwscrXjl3a53pEwD6PnavdrmZ73MU+bsSGF8nadyqjDoB+P
25cSRWPCMGRkCGSbLs2FKu+imkbA6guliW8Yo+N4EjQueroNe4lY43Gj6OmXAvAp
Rvqm6fCR3FG8G4naGH3mxv9OkfAVyrsTrY8zi/LMpN/xx7UrLyR8xau/J6jE5x0A
KWyKoarOFaimcCM0G4sB6YLBelER+ha9wlpBH6XcIIVN7nlsYjbqboYcHk0irLPy
Iyc7+3SytZDzfgTBeip//Rlbn/0j6DA9pAlHiIH018GK7EjjLCVEOEvlRZlt9125
AK3985jllqbRSQICN4sAxSYUTYn+bVkelPya0/9LceKc+YG9Jm4gwO3tdufRHBaF
B+vxzjAFcaFNf0J2JpRodXxHBS69zrmKgWVX8ZH2gH3Oz6IxZ/6Hp/ScmXaoNj1l
rqbiInbZPEP6nL5Mpi3vSrt4eU1wDedcDAVAFTnWlQb2ids02P7tlM/K5JsCsxkg
PFCRBMrEIe78ygVhTGS6yN+PX/m5GvhLspJJr00v8yE8FuPoGz54l/HPta3znkyn
/0+yJU9KSMUjrYKN4/tTZfJnhc+2RSq8VDZxPjYcvyxdbV3DX8p0FT/vlvYoGyVo
qKtFamI3a6/1n97HovDeMSt78tR95Oel4VibeyZEuCn8E+C060tFYNC2/I/iCWVl
rDgmw9ldFQCdeUa14VtwMUrGcZFfS3lGMkuiOTloDr9OQWvvcLC9s+5CLS1IZWH1
OFmMoYoR6wtQOLKO5MrGjZlxsKv+GVt61hkxPhzkXR7ZYifacJDp30JOitYuVtBy
ab1V9okfZMEifv5+D1lTYqq+JgKVOp4Gt9oXYXL4zdSlLHbciRLZ1Wt4WETQ5Cf2
OoE0B7lVS8VaNRnzmtnZ3qk1T+wHzR1/apxt195t1LV+yGw6Sjd7nhdmIl0Eiu+4
ek0SJgKM3+cTqTZl4rUk7KO7fKiT3aQJZz/5MOH3Dm43LlcYXLWkFD8fdXr5P3QC
b4/ipt55Cwx3SemIBFx5T11TLsJUme3+ljLTKwYIUnaaAmA1Frv4lRxAj7WU+/Tn
pnNPLiOUL1ExIOVvs8VS7rlGK+6Ah5X5od/jkV3NUNDokWh9r0be1yrWSDn68pGe
3ux9DYP4Kuh3zpg/LU611Bs/9NmIFRoXmU901PS7h72rtgbjLVSFWHYwr2ed+sny
eJcA+T6pbeEdAqAMXMM9XQP9CT3xXrZ/G9R/kOTe2QMOGq9GO3Od7BfkAj6BDmX0
GqjsFNPoBvfBzjOsHJK83mCn/c5RwsFHdN7e5D+abGTnmi7mm95GLdN1SMxjFyAi
MT8wXB2GB3ZatCQMusgsorgRVb1ugtvvuZ9k9oxjFfimAcy2NejgthQpMZntAV56
zGHoLk1/GH3qADM52YD0BB3Y+lgAc/sCU3DCwdzc7VlthnpfOKQ3xoPKMip/vXk7
QHhanFoZWkla/TNHUJuD4e2A4cu/gT/xn74urzdu+XcOdScqE11LHA5Y1ku+q2Kd
81dYnUV5We3E3rlTH0SWU9UctrBFM0kIKhiqZjZnWntIUf709AjNQ/JHhNxqZr8Z
Is/0mZXEjH3dZonHcHE6s/T4lwmDplfccNCTq4+PENV+EIUpwE90FCnQyOojzKFU
uYA+ajGzL+xX5Jr1dW10C4nDyfmgwdkNeJVQxJoRgqWE/jlYa6IWSdXtzNZT6Okr
Z/I8CiR6ioBjhQP6N6opaUJ705YNPbz/OLfnnF2LqFsBUsWC2GQdiSX2OJDQESFA
Z82TPz2zn3jE5mmo+VCrJ2vPNp3XektO6QJI4M8dJUWvQR3PXoTHiVNSuw3ddoU1
2lMtUWXFx8Nv52bYyYQjSGj7Z3hK+zFe6Uam7caTsDD/JlkSfP85eZfDlTkZ5GLR
neWh1mlcaOo3klQx9LWlWzPlHzUI8+AtfO/SnzUo46yuk3Qf6VMDMMUwNmVgWalg
eM5e/JOdmS9cRpKODHt5n1P0HEHBhGTFlyiVz1dwri0AlUMs3xJcRw6iQEG9TZx7
hRa6xMaXTJWATBJDXEqQsNfQAcWaDtasKUYelVlhK0hd3F/R+AKUEKKbJRilq0kY
0T3yFuB8QT0wxCU7DWSvlOYxq1TbsP7cUUtHKZ+qs0MeyPOUhkmDQ0t1UPjVS9oY
3ML9/aeEEqbe1LLmJgon+8eReOFaeVHdXhcFnMsf2zzABzpGlc4KvlMr9pdWCrqf
wRl3PpQZer4Dv/XQ+ZZsYmC79nK2x/XAGHw5QZROinVmUjFN0PQx9AriG2YNvAW1
BNAJ4NbRCvluh7ePQEy8cv2d8PemFVJZtsEOPek/+Lc1r6mEtFabcuBeBkWLMiHc
HKyMyT0W74hNJQDVYwRMYdtiVWiFnewMC2cLSMuaFF/LpIa8BZwDucpo/mWbKs6T
jP2f1fYKa5WXdQNigrQV1mHeZL9hHHkT8Z/DANiKPxaEZ1u5pm48Fp+8SoBF+xxq
kjc4R63GAXGuB9/mtNG8AG7ELwmKJumwCsBCqhEMylJu3mmAErP48s8gPwqwonMk
ObByE4aACHTweLMa0Dj4tN28tGWpl4ils3a+YX32fe6wnQt5LWqG5P90UrkBhPBT
sLOoCfPpvYPG3bgr1WUwqAMUV++KJqgr2tQm+lg5aBvO2Mr2dXEfo7ebMQjfBBni
mbwzjDBygpBmgADBpRSs1p+diDxxM4ghLStW4cE36S5I0c75InkDhDH+ERPYYbvK
BceBjXapdqKI0DvYKA2UuBa8wMXUKxrQQIEjeM9X75cEej0d4mmaPJiJyoo4ghAC
FFR0sPYRTg90KxMQNIqIa6pXxvUmaOZBlSqP27ZDfbN7avtZa5zhYxq8/6qN9rTo
zlfwecCuM6RVwHa8Ap6QxBd4MLDMyLJInUA9DsRLn7MTF2L8d1B0oBG7qiXZmEaw
Yn24BDp1zawII7yFz1W4SZTbSO7qtc5IDAKgeBNyss8y03pecZYS4B6reQ95hIie
Brrg1OEFBAeW+4qnoASiJLI+IqoO47cWYkjlOopB5uXPDNA+VUDfDz4+W0N7VzCQ
RHGJa3wx1gTlove4VSRLctvJsu64J0zQYVPOpLGzMd3Jm1CrBbdXcv2LPowVEW5h
ZSCCc1ewSGaL9r/UmU6pV6bP4+iaH0icb1mFGh+1jdU2GVigwoewW5PR+dHMwG/S
Rdt4qlQVdo0hJg+kyqIR/une6eheAFh92xwhLa8xwNZ7dUSpGYL/ny55w/ZWOE/8
wGFZvgExJ1rsuxFWxxyXY/xs9q80YPT+Mika5Wmdcc05Mp9t/Q9E+5rq9IGit6qT
YVvBQelieJZO8tGBgBTkyl5R9pELRAK7ruxCPtxjHSeJlg6dqKROpBAqqmEBWiVZ
sYVnPYKzyiBr/UNxt1eALZAPwvH9TMawM+1Mxc3C3aE3vrrmEOCcJ13gymmJQCVC
ze+fr6wqg5T234ErMrbsHO7Xm96tzJ0g7v31fyb6sjY0p4e3Nknmhw4/d6B06QXp
wPxcnN/Beg0WfOk8+sltl3PgWUGQwFadrMq+aP/ih7pWELYS6ImjLGJ5fc2GTDgU
aX0PQEwr/rq4VK+M0cOL6BWtLbkjJJWXoj5a6fdOzC8LcOv42Cc4h8KgP4RNMNwy
nZhsDMJm3qQzkAZGneZvp4FPtwBx49K0LiMZzyc+Eo180n4RYiOQdZzxvE+UPd3d
THjJ+9tsMcaS3+lOw46I+fFLlXt0iGi/ppY6vXP/rdh0PzOwNi3tXUiOj1iyC7Cd
ACCfuJIJ5wfgEzP3FDMkVHqfXh29LuUyIs3v+e6Tw+TEBHgKjRix5AK38kxMMlqb
mfC7+TSYV0hbZDijO2Wh1jEQnyC6IhP/4Bd5Qz6EE+MbXHrj/sQVCfy1A4jRQdAh
8XzOYmWldJN3lNTBUtGZTNoZEEyj5HtgYEQnggKWRgwHKdYek7py6fSMFg7L2d1d
5cDEbG3swnQpMDIUqHgu0dNtg5O++nxawhzUZYeXGracGFwl7K8jvGBW72lMd+vL
ubaNkv70ncIkyXvqUuStt7OA7sgmYWl5s9gvVYChJe5LluuHX3egWJ6BY6zqSk70
C/hF0419uuf+e3FclGnmRQzaV578UFYkOQZLArAFKMElukpFR/ydU1dGSEl6nlIy
lGWkr+EuWW+wmQXH2L9JxXjALpKf6T0sOcuSXnlSInbqvVhslO38232h/Qye1lav
Q/hxW3s/up9fDU3PZg/7jFfoL2DvKR09La/vQysxa7eWzk/SWkXmZ137ZP/uiFQ/
ZeBJYl92qTuUOBHhVUmBWvVCgye1rf8r/AE0sDFpd7yHKirTVhzkjmafFIQEjsF1
oq/OJ5PBBO6FoC3V607enMAAdZXh1+HWGbYgGIuvoKeHGVkoSayFNqjoKvmTYIj/
KKkWrihgxaZmJDuf3n8F3/JxS53n1x8ed8mxkxL+kSydtnerCWjLoIgpuR69Ucta
Pkqev9zUdKdNUnPXlhydmmb5XTdU9O39th4qhucuLy3dDfFcm7uexgByBeHVclpY
/9qufMUsCqpYMZ6uhdrVVjGVC2CdWXb7zCuD9X63/LjIpGdiqG7uimQTTBAhA6Va
eWW7HPETjx3SDJ0WiVlvTGcQpMuIqRnOBjPtuekb4/UlEg06OHGg+aGYVs09zRgu
IFyUTS/8Kx2TpJ1oZIA9KzxDiIzgrmyUQuVM3xatXwm4TUVo0S4Up+bcK97INjFt
juYd4k9fmj2wS6p1uh2bsGZgDgLOw4Gu7yHmwDC0mY/CNXUZSE4sYTPTyAdCScP0
FbVVXEUXieQgTt7uFEB0HkDw7CXI6NSTz0gc5OrrwOKiDhP4tOwxE1KH3TkaOsz7
HiFvuJf1EP2e21VDsGBVFF6SNWDFMmFVusDtRv+X78KZRhBOWOyLTdaB/4RMEQsw
HHee7aIyJmVI8x53dct5yc7NGRFfF0NLH0EFly0Ufk3AWPr0d3UBJO3EVmbMHn/Y
9uIrfWUNQTmC1SM5otnLm742GsEJ3M9a8BUKnMHDSeWVBk/6bpDrqx1kjbZwiLng
h/ANs9Tug7jfPKpQckUvgj6MILWfWEVS6+xUuMLpi8zk2JibQZ8fVwNnx7owLaWA
B5BnyNRryyvNTpX0HALktWuBuc8veyFWcgbtZl5KNro977QsCs4TZsfYqeg+Wl0d
LWfT/FnQoYRT/z4jOym0ofkM0AFwEPGEim/5wWNTUEySOV5/7224JFi8xBLhFXkp
LMgOMmEEwUPpuS/J4Cpey12URXQQJv3WSZLNvo6yiJYE4UoBrMQkRJKUXZrGFXB3
Adtl2X3Tj0GNcN36uuIa2C080hInQ+13OzggCyKdar9xMzG5LN8GgDxe7wSDGU+K
OlUe2+k0M4sEB/0Qzx8DK5gWYTjHaMY6gleFe1T1JuATW5ZqpY4TLMPid9C+Dg5r
8hWA9uEWYo5ucanCHYS4Sc6t2fxpc/YtvDWQNlE/vMXbJtRXoM3FNV9d6ydlJO17
Gp3M2uERFuzJZnJSA5G4Qioz7ix0pmcL0/xBq4/ZiLOxjmAxT9qPWqSxEu5dmpI8
yxtxXrpnbMVZqBZrnMO6S2fRq5qrH/om2p9Vy9t9ACN3BaffUWENUKsNnRWS5DFd
DH3pXiKwumjYYJg0KWc//c9178PtqjYo85c5XzMfhEGk713FA70bN8oMz1SwKoZB
3glx7o2ogU/S+pwwhrG6ZLh48iRlqN5yIbrJf4pzC3L6OWQGYD2J4jMtivCIWavZ
WXmCHdT6mwBkfIECHy66DR06IodgnJA6eYIjAttX/d77xIgj+GGbEtpiGie2D6BU
ZlrDdhJ8ymQRFoDDaalaxoVzuw6O6kALNMe1eAyWm1Nn3In1Cf5zW4pb6fjnpCQd
KplHFD63hSVTxYLPeyBri7YvLHVU9SUNALqUtRyW5no9g7SZ3fa6SkMVqLKhJ8dg
JAh2FOdL/az1B7jZDVhB9NSvys9GSE31kWEUQlAh3iSy7VvU01U/WUzVB9m64KcU
hf9Xt9Jp33cIlGUauqseDZ1KgEpxsdVUrh/yR27qaq+56oBGBrMaIelol2LMlhim
Lt1wc2zys8p9a5e1EOpyNx0zv6rMkeMVPsJensnQgQnseF9flo6DqlpE63Z/vIur
gwrO5KlkxXn6aPQZonx9NZZsAyI1VlxODQyFdDsdht9hmiCZnfaJ3EJ1eEGXOXOd
I/4EcTFiJ32VTLko/F/iBODu+hsRB8QbnxWJWUfqI1sss3gmozvFL/rjbRbygTIK
8E10pW0QZ5eJDaBLv5fkcUpnjfS0AEEm2xB0Tj0zQnSDjVNEFZ1QIUrXGKmHAiwS
WQoAvFmv/2OIuWiaHHSS6aw4awrqWAkTj3EpxDZPiCmscSJkGinAyz6YzzY1v1mY
h6ZmlBake9JUCWlq8hrkhPgYYHl9kbEkLfXp7GQsCTl1bLGhTcs+eo/fVEugxL1d
IaB9QvU2o2/80qFOItrSuYx4Vnu86hxf9SIxyLurOfU3FL6crrzV6KJVYyKAglI+
g5DCMDV4HvsyERhBs6If6flwSi96onuMQ9jmFb7uKqRqw9hKLcPExoX1iMQje963
QWN+ZGnay5YwhSt//qv2jJsdvcI5niIRzxYcoOFvSqmTTbxxBbbSEtl8qMkac5g0
Hk6fjGox3LWUcuG2aTesaCNLS4ZVUvF5ZTjS1cfRtxL2wR5/BT/XBTX3QBRLWmGE
eIDBouArSZ130LBmib6NL6RIGIh4Gh6cYHbZpXqJ+LFt5tGE9IlN9sCZLhUN6rEb
+Gy02cEF+zDjy6MM518cgBvPFvIW89X/WMgpwKL66rThLH8hOjb3uxOgMxlnfgCf
0zdDQ5X5jA2cIbVPdf8OHVqdqJMlFpCDbvS68+Ju9R2WDJt2DRcf7+SpgANvEQVY
pGyOH8bnYXTjx3J72R7op7uoLFAvUxKYJ8yvOjkYmYHsbg/kXI0KvHbk+v7dn6g8
HzpBATZCHAftAweQFw9JAZ9JmFp39nYN2lz7HuDmPlCFihnFmGEVL4yQGrRzcmDw
Gu9QNJefYm2AeIm1mwk1cQIeht1kK8i/bBC1U8u/+HCUkXVp9nNE7FE3Gy5wwsg7
EbUeduRyNz2Lgbfk0siBRje9LuD69pELkXpEfK3R//lSLFfKN5u7h9140a9rIsJ2
Nojb5LvTZwN9gR+D6DlAbEbmhD0VN0WzA36/csCbK0thus/braiE11w5tIljG9jp
97XcmdNLjToEh6A7zWt2Ka4pH29/tyo3cPyqRyM34baS8VGqSiTxJcnHuP2/WBkb
Qo8LlQvyK7XYRDpQeS4oNSAehZ7KRCHX0y9S/T4pub6x363Zoqd1MyYvVw6Jyo97
CneaBGlCanJkHPPWvSkYwgVH5vGOSBy/BceVwifVqYCfEO7jA8lWnzdzVehHf1+n
D/+3Gs1lvaM6HMPKZB+IYMSajAhszDkdelDSLjfp4JlRQiIVrdn2RZZz12C16iLw
3Yz42J39TPtoPUx8XfJB50sRQxfFDOHJ9Bb0RCX0ycMWxw/GRukktO+o6DmhjOFj
W8baQR2sQKFbEWzlMD3fu6f19lPONFUrVPqPkmBL5VaQYPwxEBG2lOjhLtRgSD+q
TgN4Gb2KtXwFye8l7XmmfBGLyHwBahersW6YyRWPHh33gPdBJt4AP6zuusfCLr3z
nSWfxw4CoUQ413o2eWc1g55Skr8rgptbzc/bsaFy2/xSQiByhvABJoEacqelp0Kl
oTC8VCB8zCo/8T/7sfNJ50VU11I0S5NY9dCfl89Pc24w0dno/Dm+UcV2u13+gpIJ
5g9JekVFCXW1/d4jWrOsaHW9o8aA0CA2Gheb+GsvvDB1Fjy36rMZKfWrykAdFPxs
AawC4oJH2F2Sfm4nvA8FmrMXUsxpb2TuCl2aBd0HsHLAjKGWdmNNVi8KA6VC6s4e
nDgVGln0uRtsN9b0qMX80NbokHoXPJoEKTdkTKMXyu4d+A9fVvMjnIOXQu+lh+n0
C2exiRBHJfuO0LVFQUeYMles0ram7pGvueYPcugbL52ht/4PoJ0FlWORHzKrNZhR
aOfmhWrSUL5m367xpWjzkjtZdb3+hml8nQgk5mYcY09keWF8F+ZJkwcn2Ld6iWBa
WgHlWF34yLC9OGeYQeFBJTo+k1THRDdgUtqngjhXFB3sxqz/Nc4zJ/uSznImcjfH
etYhbZCJ+GjbW3eQo3pBeWZuwM5GbE1/Q+00o9MD0nUqNc+CS+ANCgl/TFvVQqxM
iu4dF+GgtM3xpAqhYWZsmqo/6C0fKOhwWbNE9zn+zOR2+XWNlMpnqm1MN1P7DRZs
y658nVb2S29mp0Fxat519ReOX57B248u0LX3lf4is2w11c8i0ksSyRpzZBCcq9hx
W5GUg5CwtpJXRe3E12Sfh3HBmzgQ2uNtV4DqQUA3N1o6OUNmmYwIENUtxcQd4vse
v8Y4Xmdcr9Fi2lQtmvFyKtSYOZqE2Bi0B0hFTmwCHdEPma1wa63AXBHgiKbBos3r
+h+vpGTzN5puoVQaEh8pOwf26j6ycQh/741ZhUo3qgs1egc26QktuIS/6U3gH8Xj
rVSPMpJcdDyaahTmQKfQmCbCAs8V1tbgINQ6QDmpXwISHi8zRdHk6s72TisVrw/m
ExV9vG9A6rBdRrmf8OektiXFga0miPrX+xl3cUlpj1P0Y6wlj+PHvBYSsGvc4fyK
IiUe2dWpoAM3HtMPE96nu/lXq88QewK4RlbGpHmTc2GubcHml6cbj3rY1nRcRsFX
ML62zUlsOqRaZWAahcRW9M+Kjlk6SyZwNnxw2U/f5dD7KITOBWepEytQtjBajNue
vw2jWBYsYsRm/ps1DezlgGb7zL3VOO8ufO7sRyvM/E7Zr47V+waerCDiv0BaYLxB
NqUcvb+gsewkP6PFNnnFaujoeXDMB8KQ2d/9Wq7TCmetBXeG37JaLXpTdpLHSg4p
FHXVSXS2qhQpLvNYiuQ7HTF+Eth+WxzU/hGXQyCWSWvKzWYKd6oKAUo5UflDp/5z
wdGHNaQ/Vi9/vUJ65BR2UGx40Bk/lmDisHbyCCIlD/RQhmhOSqtr6sDNd/nBMUI6
Nt6TnN+RxgH3b0eFQyjjE8pf4QhUEJBA3YRwBEDKh1vlo8VQn5A35ObKeyixFBF6
SdkT+nBFXtuzt0d4ku1TftgwX+Z5NNyDt8ONRpYQylVqxjmzCh/L5C1Af4fbbFDy
m/9UgzK1QdLUMmJsXbC8Nuc7HLtBEHiHiopJqoX0RvUGnf6+I6mDwXLSjsNr1W3d
PdbSU9L2wfootgP2MeQ2HBgsyVdmaJ8Ew/DfVQXdLakiV7sBXt0sBiYqx2QYiazt
o9WMQN6/TTUpkFYBAS2sr+v+/xQHHHGHnGm0AgLNK7x+a6x80YK1zsPFM4gimMUP
h1lj35tVE3RiHxRIeKjYughVy2GYsf8mgZtT78TRyPpUdDzg+KrpBWO4oIrc/083
OhFCls/wyM/BuKoS497WplDMkvSzrorZYivJKlYPfn2xho88tMx4jfbJrwlh83M6
AzcBmMVTQyWKIAdQCzHqHUQfA5BWC6IaTpv0hPg1dUmWfk6rEW5+sv0HW4QfGldy
uJjIsmJiOIu1WaGLkX7P/BJaS9nqeBCdVcTZN0EtZivyBbk4Q/ZxKSwpwzeI5ThC
3LhmbW9O9/RCv7nHjvXI6KlpCocaNhOb1SWgBWglVYvBfNqpBGCsySgUpHLwIbTD
5M7LO3/ObbMzRK4702TwQHr28g1+J9O0XYvkSlmEsMWogfvjdE7VYoEPk4dLMFOR
ddeUTAMjSZRu5GeztTJcJP3XXBQn5ObLROyzCgLF4MRkPnFED7Q3L4yj+pDfmLTm
em5IXl2GzDTZ6CHhNFlrXsjH+zl8l+dEIGkcDtk2lqifPAYgkSoViQQLPkptK/cz
vYPD9JVOQ6cywGWCEJp6DlORp4+Ja1i5JmxqCkFM0kZdpXbO41lxX/zDod9N8RBW
svbI2Mw++VRItkudeH9Dc0TrVHGnKetf5LeSwlgv1ho7+ijQ4TN3Ke5qmt6kltBc
C3RrRpwToRkoOItS/orBfAadJ7wOfpLbbOpe1Lt7Qv0QmmV88buZqFX3LCHdD21i
yRS/yH4+SmC+iSlYsexKhJjurWwS4M/8eMgl46RxAegsLpawj6nxSZ+V4R05O6Uk
m8qgyeMYo8qkGgcnXwS1MSuO5Sup9F2Pe7QVgfskufDT3iXUFD9Uf4g+kvILlX7Y
GxbX3gMqfMkYArSN5IlD6ofimGbkiykov4eO2u54hqpkKe42UAq3B/KvTNkzn40c
4LIxTF0uwR51wuhzY6QerWKG58IaHK+rFjd++a03ykC+ND0fGwBMPHnDM093LC2D
6TMlcTjDTI6xBie4ninZch519whR8GZCHfO+lN9MhslCHKiOn0mDubly5PsMuiBV
gC8ucrRxrBtMDPl41YauCociNTd5m/5QdBkzFXLISp6iNdASGXU/3MEdk+AX61xk
7SAPdVchwRjsmCIlE91VYaibc0V+ws4rGGrqF+EUiq/pg/qlUx4KsuQh4XPrmTMD
3XNEE5mEXjciAZ4vMBuQdc7sjjC/vNT4oUY4tUu+Za5ipwLo60kNIwtxQO8fxlZ1
VpvzCxtYmdEL6IazSwwUqWTDVGrOpNROCKNZGAajETFVTdvFfxHRh8p8an0inUhU
+eIryG0vGsyKCJROXmj6J05UmV2wJ7rCObuCxOJRFz812kliT/9gHCErvQXJNPo4
Jfque99pzPh0vkI1PGPfyC6l+dJv90AGZ5vi83HSYjGNuzFZEMCnTLgSAwsZTRCy
+s0GG51R8TRVRudtTpTtDHp+M0rT0Vj/zmRc1mxQYQf5Hdc57ebZKite8huPNXUs
4zITQxbQ1UielRh1KP0ed0gM0dtD4kLD1dWpM7b2bWP08DamfnxO/l1gpxPHkNqx
xpBoKQmW7NOFLR4zND0+i+sLcSsTKQqHalfchcRoxQ3I1pfb5iHP4j7xCJOJ8V5m
9n16euWXfp/yTj8ZHyhAlFIB6A8aQCDq1hDx17T8fgQZo7ctemTmxYNs4vFPuPWJ
xSbD3dbWLKJ2g9YwKB+vKq+ScNVpUYGEpmYef4xds1vfHljlPTYS5onDHe1wr02p
kevfNCM+d2Qued1pJQ5gD4lX430ROwyjbQRu4DAmiu8+Ghd9bJOtVXFZp5mlD8Gt
d3yscOzsthLAQzeKyCceA2sbgDb+BfRtPZtmrMVvS3FIUklGM0zOEQQGebh+QRz9
RW+r1aDc5yW02coYTUlemlsADIBemRJ37HUWVwR5kpqu+qX+qDMPEVlgR3IG1NxL
jL7WHM3J67dmy/bXU9I92YqLtypdwkdEj8r33Xx9gAi1SAZPMCNUNFf7oKNsiBgo
ygC1y36w+2rQKMMbQ4Zs2HuIB01PUfsM8p/n6NTDx1OWeQb8v+A1U0PpT3ollVwe
g3tn2L3aU78cG1agU8ndNIXR9Xea05b4GYshw9Frf/O0lI2trStYaOHZ7HMecjW4
/rdG6fLV5NTLyYp7sSnP0P35cuWZB2g0NSOlNEMVS3lpJKxvQn1UfJbEfOHaxkJ+
6MzTP8B54ySYd147oGLid1IhTMKceKX25FCe+v9TXD5B/ylHQKR30GuuVmcvhybg
TtrzyK3qsUOActFp7eyWGMratvw+yrndYhGHCT2Fa51QNwPnMj/07R4LjC7sohQ0
NHNhUZ/k2AR/jEagii9Qf77f1ZoYy/FWf+tqaf3Eb79LrTTwGexWRRJ4e319sDa1
Yk6Y6Ik1/GzZFc+0ggHE0iN96q3fKIObVvKF25NpuPZkQGRqwqxxWqfkiz6lZGlQ
0sQejqP/TopINapTaqibqvNhqdUgbdoh1y1M8QBXmI+I+1Tu4TSH6S0VOa7eZSzW
26l75Ry7PL5e84zqsvjhKngUqpuPf6jUbWHB14SqyDGTHRj05kg4hx/D3z4loFk3
0ZG6FpRpzRhMRuBMPtKjXDz/0yg+raXysJ2cvUC+6q+RV0S7Zog8+uG9sQaI4dr8
6hYoSO8sZEHyeSgMgeJCH8zkNvxioWitFeHp8nc7Zsy2b7vfKHurxi8T/ntM6fwI
klZq7HzzYGa7xk2ky12Sh3g250F18GNg2MihXUKNTsczkWdNDM16wXh6LPZ11YfU
2pq+4Z9uCqpF4PlSnpGbE4tZzWTDT+AuCLLlnt2Zc3JvBZAapz/KOpZRL21bza03
L44iUUFLOSUt6PESDVBQ9idODCsSeIx6nQfImSPb+3e2X7eOvlUySE9zGMDqO6yr
5xTo2SBsD96I22joL0M7L79Iaz4yXFe4NfncZkNJaTBduTVFP2iCMYPJbv5edA3u
wk2sltkC21GOWZkt4S4WvWlPvuYejJslbbkloV5wHfyF0GxWtBkIrI7ChbXGK5Ra
0XDDbcj92RD/cNhu3aBghd39K+tLwz7SRjmBvQoFh+ImQh6uJwlhlyIeIAdXbUbU
M9wFqQ5F55KBKWoFDeZ+zZ9JcjWRXM+ei6va/Gyku4M0OmPkUvvqm33v78wsiqib
ys7rWXzvRlw20Q+UkNAef8Os/jdSXrOJOF3BRnGjQ4ZXMTPBp/3Av5eGWKYhU+D+
1dJMnpHc+izc/D9/sUs1ptk4bNISr2crhVgg7GvGbIJBoAyNj3ji533taBK2utqD
QBomedhjVWr9h5BLwhoZMOILjSf1S9QuyCcPqNr2veezbm/uFcpb2Rq5JtDw4Hmm
Sapnc15h0hOnQ1MKUF8SDQUlZLTGj3TzWF2Kb4NbpoTRzhPRC8gnMKbZ08BuRbzB
3Lk1gBKI36paBrPu3EoaZjCQmmUxg9fLM9MhaUVhqJvcqi5d4Ntjkzc19N7NivGd
FAPqJTicKB2AmJvm4Yrt1IurzQweQcv+J7a1VV63CGg/oOqamAZIH0K3s/p5RFj3
r6SVtVVSVYA1BYCBWip4Zunq2kzd5+K2lnZ8QkNt35909rzkniJVRcazBgjpqFdS
/PivGlm6fn+Tw0TLGbFqm2p38Lyl7XdQ0cN7Z3lKESxKxf668/Sxb10quXX1Ks/2
ybOwglDwmPxJnQah52b7bLyCJBfvoUflF4HrePUBFC8J4ZJaMikAp618Zbpdq0Rx
2FGSa4m7FxeozhTmSsZbFLHRERfKcxEWMm83aW4yXdFk7unU7AHDH6XJpi8tLwZ5
HZGbvVxMiLOCDWRSSOg/oRDRnHzzLPqVt1caWPsZVCHiWok3Qa9bM/1Lbld6KNyC
Qh5cA/vT5ONixyNtz+q2fNDhl/+a2n27CKsjxxLJmRuNCa1db52JyMvnPRn988QY
dhjpaqsOFApOtp9Dgd18uwaVo/3qW9KIiSVef5vRtQ2q/uj+KKRfz0GvBAPuv5/+
z1S8CKr8tMkybXcezwzs92hYRskoyamz19guUoHrZJtXEOB743KNF/gQ0DK+Vs+r
YZ/Ya8yMGpQh0NmgE5Rli0NWK5eTdOriOQCvWFcOE+MOqBNQ8wAq4Y7L75tR6VIj
cpAFJPVLpLggf3mpaX/Ah0aGMTvzNKUQLSWeWxrMXIyEq0ZG8kxkMZsDVf9ik7qq
G0rbx2jq3uYBX9IMpCKXxQVxoWh0Wb9nH5/IaqMJ/jEcGA23SWMtqdMN4U+QaE/O
kRJm+KxI8dnHfQv/5jV63Q9BQSph9/tB3noTe5O+m3ZpngezznycrItTJTKxalT0
ZPU7Notn1/qzn6R1KSKhTD99bYPjSibKmCWdChwZCk0BOR9Zd+3RT7amuw8tLwnn
BpV7LQtu1TXzJv5koI8q0zZs4zKzueEjYyyJW9GGqI8uQjfYeT2Fy155OJ30nzmX
JE84mAmp5uYy17JveDDVwX2798R/EwcZVE8zPgoJOgGq0bR24z+k2L0lYWqOabqG
kdvU3u0jefkrA21DEcHGONw6qx9Plep+l1wzyezfStEdag4fVZRPwbVzfZKE2uRo
aj9Oq3zJIG3cf0XdWN1Nr1/Jzx4mIi3x653YsXBxpACV68AGl4CzaFWQLXQKT5+z
70Y33j1/88wZrrdlcM2uZtETlO6Mn7hKedlvDlr2njZfK8PNP9CqcUAGjlxqiO+0
SpNSFca+K216ag6K4jsdlupHS5i66h+MKshY1sdei9rsuhXQO65gUL/pPlie2aB7
WCfA6XgW+9JZByR2RYzEfAtLfeDQPBvJoUFrUGz2jwE0ncsiQD+OnsM8ZpGv/zMI
NzNM8QCawG1E960o+ZVYRZGrus1BIT9Nkrs3TURINNqF3qSgQKDaLtW8/02RVp39
uwnqDq6kDX8FATor79QrreblPzDjSIfA8Di/USmw92q/Ajfnxxy0YAohzKKAOL0d
eVrL4DOzfGmynEJc0K6iMfIxRkoMMGmVsqOyV+s6f3+Kudx+dEuVIdoR++htAGxg
52MLpa2e4DwRPFGfZcML+BPflaZkolUZX3U98fbEDoffXRiKyvRCW6bnnLCPguen
6zTBZSxy3iBFQiQjNFDXNCEcMJsi475sUIeCd20tlu8vHFKUEsb1px9ZKgsRa4M8
BmOuqLYZUPRDj4S68zHSEg7I77MkqYIB+AbgT39GOTUsYdpQuARtyihy+h4bGvyw
GaYVERBoD2LI7fghTi8AzK+6KZUdSegbi13nDdGa6JjFno5gOY6vDo/yTeyHDaOt
4wFY30tvRCkzJmkgSp8PrVoCuTYkNjM253rJTykQhOVepGUHmmkZontc3ldSrBam
v6mdpi1IPrSz/PpI4xXFGCtGsoCmG5oH4vMSMf1g9IsCc0NYPWSfQ+iwEd2SDWs0
kiRnvyH9zJd7A20f4GfVvlb6Y7JiY1jTMlc33VFA1IfHOJp15fP8U7k4OtHB2iWm
4fmULUvljbPX/7PUfqpGm9BNED2OL1ln+v/B2lm5fzFVtWuwTHG2p5A2MxtunzEX
McwNH9fxw9kZeNmXwxY2g5mKSxZ66BlcD3jpCAcrbhnSt/uFiu9NPn0c6NHEqm0I
OUpSqGRo+feqU43OyRB5OApxPx07//H48d/TRxbcQwJrwH6UVR4rt5g+ASFsrMuS
Wk+KZC0YCjWydyRw2cLSeOb6vpblvdn5VJh18YF4YOqOxTExU64Kjd2C6RsTMTjf
NP+H4kzOoViTkuzVj7OxIeoXHQQ7LkXUJt5MyV7kt0RP7GJJg3tdfLRGkGGtlltk
nEtyytEHnbZIoWlYvIqRBjorrViNSagJhU910KSb0AkyRItvgNImhnoZE23fF44X
ORitVAxBonIL6k/Y/3zk3bWm5zQSyqRWfLdLp6+HX9Roo6bcox5vHFXD6q3MWrLE
zNmzuVesDteet8vkhs1mdvB5kKxiQVG1cK2j5LUdQaZEljYH9EUap60xzH5WE1HR
DMdB08X/3u3FYIFFKRquUhJRmEu3tA1ic1U2WVw+dRl91MOhDFNZru77lJwrsHIc
4mNckfvUUqUnoHMmgOABK7jCIe1bBJBUxYkcvIJRzdb0y6n0j4eOLCDKdYWo/iVb
2yWksGuPzD+puyFJmImNUqIxG5q0A/mJzBbtvDM+aSxWf01kASYPYV7BOdJAiNPg
8Ry1DBjegRWzo5wF8ZcZGyrDSaEIXB6IXHi6wDCZW+nVTqRQxU0u/P+AT348/wLS
M9dmPdI2i0VpIGMNjqOA3Uz0vcJm7tGEjUZ1ewKE3c7JCg/W7W+1YSBtOEIoAMxB
eOj7bTsIw71p/EilWCxf7GbY2KEVrZJdU5vHoUdKnJbFLX8R6+qJ1rX1EcXYe5XN
mdiLdI32SD1gRdVYQu4wTu0NnvQtpl9mE8lNhWcGvnvPr5YPLQQ+T0eNTHIqf2R3
xn/Byr8OCpIbWyuIUYv9r8WmY1m72F2Wp7AAuFOEJs5aq8/19E/9qYKg555bsWMc
Lx2ic7N/jwJ/Mq029QipcKL10OND+eWEOoIvt0x3BhAkRNKXNwq9EihJIti6xsDa
v/uLTL32/glVxII5y89oDLSc0ZbjoZgB1bdAKS1u0xjXsIsB8QNQuGGHTIHdKcmn
N7fAZ2uTmIHprm9fdZBeIDTqWunBQTZZC9IRdkww/zYx/+WR+xuMXVxWWJ8HaBGr
vkJMvUEEoN6UmQi659Cy5mZfdnbm3sx1i/4+BM4LmNMTm2FvhG9JBMO0FIHbCv1w
7nguNVcMxy3jLtjri/hhOQw1r+PQc2yI9bsGzCf/+k0WWDHUeZihDIKh56mcNQ4O
OO5ILkYkj9trFSq9ilGKDEUUusHVtky3DqvFZuLqoWN5qHUzPab+FkUs30DjX4Yw
xjofVow1hj/T3mVz8qPSJ+R+bpCpz0eO3YT5DEpZpBaf6f94L+L29NYZlc5DYZTo
9magq/7ZazIQRTEG0F7jdYZK78H0v+4tnxFWoYtjmc0UAy93b1Q7jDw/5TSqHcFL
/yJA7u+CYcdZVqDeJEnkYk7C8p/AiOiRy7HEdxyZydA8NLp67XdVzfyLs4WSEZeZ
HMKRzqdszJ6qh1u6+LRvlWnDDot0LE23znriq8hRAc92TIqS1O4Wu6BN37gxC75y
RSeHMPOvJXk4BFUIpKUlQ5QLrZckJ7sckgyKLrm+taCS7lq55Fc1Wss/VjZC4TYS
uFB2fKA4/LcERMkAfZsguYuSO7sGUWNqUlnNRjDkgfh7XfYGqBCTOMlp/CUO3xGL
PuAzO7tRLuR9Cyq3rw4ijGAlHZ7hmY3ge6ynDiWWgY/0ps9QjHKVBYGlpDky+TZP
UAbKZcrSiUxEHUVtPOVa+8qI+6sekVsVcWvSQHgnm8ed/VL7+eKuW2I3Z78cco6T
or56ecF7RxxdqABtmrpF6YT5wqC8dg6mFy4RuVWvXfucGBUIIh6/K8R0GBSfFc5/
aIEIW8iS/tI+D49NiKLn4qmpOjs/pTlvDUxIO1P2C0E0QEz+TocODBuvxfUt/QUN
2lpU7GdzA3MMrXGpPGYqWe0Fs6YuZcXE5AX9L06EnStkMa82v86gKO5oRFNNWCBT
M8tRF9ckdiapFpjB+vejeBZt4/WHGpINb55b/dUQnoZG6+1z2CmzD5C/opIf+K4i
kyoWUVASM04s5hjDebLSuiDKTt4Bf39b1FIvw0eh6HJEPwUcZopzrsj0UC+6c5E7
gzZYHsJ1wTxaTQDsUVaRDP3Uz/NrDNqeSZ0mRJPpuKK4OKd1qk8obNB7ANN2Oqnv
lTTwDdQ51apfE+UBO85ReQN1cKa381veTWB3O/ZECFoeLN7zHrST2RcrUcSZxbbx
5b/YwKjKosmssoMqhrMmqoOQoylHMw+rm61VY8o0s6XK/JGKndLzpw7SoIn3IqyI
lTaWJZv3auC7ZjhcPBslq3baPbB8xdzk5MQ77AsvPa+BiEVl5gpsPN07iiadcwJ/
YIIbJ3BitGTcgH5lk8RgV4uqDom4wLZssuJ6/agbiWPc0GUDw0o8jcx2vKx/AWAk
hLWwQHqdD2pyx43rhtBoXP53i40zaM8BuRZCPgqTP0cs/rcUP/NKOCaFLPQZCbwh
uHYnWAE7VmTKi5XEmAKLG5Rb2TMqbSMeGoiLYWQTtELs9uIgT9UZzD2LQGfgCnd4
K7O4ByeIMhkyzu9aaqpNyXpQjou1jO0HCe3OG4i0c8MTCynIm9MfdyD0H+ahvnLR
AFTGbqGKKssaxDINJi6CNuPlDmHFZmlmcQKmiGxrk04G85XBwKQqzCEXsttVWzti
X0jv7PeLcafRmzCxMNx1RUyBToon52/DbDRNNOZSDlVYjD6geG9jV9kBvlxUVHA5
ju5joeU597xzwAVi1LMgZFsQoCko4YOC61yNmtdNbVVeN0LN7YZdi1a7grX5fI7q
lfQ0jJM6nA7uoHbmndeDfYNO1d1ukiuzXnJ4e1s05UKBV6wtK7uqsqMWDp7JaMVw
0jvUHWLunIZBybS/tx3Ur+LHDIoQj8bqbK+0WpTG+TDqyRsEKiWstuup5aSSuuL4
1KWWJQhR367BrFptxKPsWExoOJ4Z864GaqNS8ZBiBru6sRUbn36YiyCAx06ktNkE
Ou/MqqiRAyLF7jL1hD3k9whxp4zooM1IUenwGnmTX8te18uNV2u+zqLnMlMV1axE
KnXE09tqc0mlEuZ7pWPWChl5gvdSgedlkMB1S11tqo/xlBr+Jk2S96sy6ThqXcrv
++HaAqo4amcflmHefVbe4BVLVCm6Qqi4CZhwYJml45zmLpiFT9IhlffrNiwV0U4O
Eh8abn8UDzccN9Dd6rCht43Iqbg1KfpPM5KLK5pSiCyPbpPlJNqJWppp1MPPLIG4
BwxUwMOI8Bac6xRhgySwNa0h8U3flOo54UtonnCxlHhZWyyZ5yYJNURxsyhvYqXU
rMBc6/QX2nePZY7dg6olP7n4eTH11CHMEOGSTf+cj9k8J8C509r3SZxWsGehTvjw
/exX6GdG0A/8WchcI/3HyGF1xhkdzAGa9xW3+Hm5bUu7QWEOd3e+TrDzeZH8ZYUT
gR+2zUXWyrK3r5OPI+u5fZKPTfZfd2X0eT+B5rnX8hdUtWbDDCimxp/8aFR9oCKF
Wenl535Uthw9/gldgwpTiNzWJWWtRl4HJ2n0HY/8R2ypp4FgufDcPIkeHjI5JVAa
4qkAs+EVBBkJV+GBWUw8E1OdMj1iWw+UkcYlh+P4av8z/GoXbTH2fMOp+GBXOhvU
dRvI8AhhmtdKkBMr2SvPQ2wsgm03oKXvvpyadCJv7QiZG0kQtPtn87Id1qAxCyEC
mQ+vklGhmYwSL5qTGYV4FTqVnhOobRD9lFWX4d0WeC+VePbdtvgRoE4qrAs7i2J9
C347KzRM3c/NhM1CySX4Y0nfUBqDHpV4ScwP6uhcIc8qh/DujylxyM2Ztpd8shx0
XGhhgNcLCi+NOI3vxZcBc4MJ7tnX0YSCxKYdIkieqStvqWGf84P4XO0Oir5qA9mi
v5DJddpkPM/M4ygzemVtROJk9DRvycjVeMW+zvm9ZpcyTiCkDX1Q3p7Hi47HsCgO
oJQMQc0Y6PJYZqVA+8dspliuJmoY0HrGVJaHULXFW9NlOM2ZRWzOweLjROXjstkE
WA9WEx+MBopsx7N0W/52W+LPwteNzJv/HtdXDAoaFnoX6MSrIn5MokW09hjYroI1
0CBESMoEspa/pWFHKyMXf52UWAtfNVZSJNLT+ahSQgrePyUNMCVGURMT8FJXOcTk
PIuWqJhpaoC9EINXUpLXzBsXnqa9T8TPNgtlEi09bo5oAo6lt0L6NDiTrr5w+4H1
oiZKIi26PykVx7a+3v4sUXqdg211Y3ZBTKnKi+P+nkW4PXjFbddoK9sYKqA07PpK
R8JA7a72evFKIJnO/xIob1vR/2bb+Crp+N0b2cJs/2CZC1FchSgUAUvQmWZ63+3E
w84J2HJqt2VdMBqk4PfP5K3e/d5kpzoNNl6D6cOvU9tXS/kDiywCvqtJbU29IiVa
twrnVNZI/wuMv/f38maSt9AkfO1EWKzOkKEuJqKkkh3iGDLVVhTp8SphAL8EbGyn
Z81H+RBCXSQz5qLxUjIMSdWxxYdK05bOJUptg6kt3AvXwMEpsGQctjHiUi61p90v
lgyaiJ98Xc3vLS3bOwVNmX1GAD6Xu+DHErIhoV73Sv5vq3/JnwWjp5jyvsVXqyXf
ZNShOrsofgbkMRVaOVGOdB5ZG+WZlz/BKomexqdJLkf/g2DzRr/CyY2UjDfVHm9i
G6NHVxhA2fKgmeImSqzWsor9K5VzGyjiBSDGpgNun2o3Q027dl3baCBRLedUpJVe
kTXcpKcFcJ3sgxroNMUZvjogQb8GJeLXWCsPedn4aeZYzXbemI5flH4ZIivkD8gQ
LQbALweqiUCMOy7nZzEoUXwZZJCe2kkWP8feO00QZv6Wi2ASM0QltopoZhOQ5lAI
M+lihMh68AcrX4LM50oE6yYqJlH7pEaF0YMQge9MzRDZny8WSao2G1as8DY8x8rW
JH++pbrlKkbGFpBq9VEbmNQjz2CEMN2lscvR+ici4FB+Wsy7bQKyzH6a74KoO0dL
tdgdm9oWbBLn3qPhPkyQvL+sE1Roe3eOFDM/UWlSyIxZzU4frGDhAT6dvC4Peq3b
shtBkDLIY54y3hVtgGGRP9TXe+JS1edyEiG1gC4RZPk3AESohkEjSLRg/O2g9be4
P56HlSoXyIUtAT9eMtjSt848FKTSa5RJpPZ/hszIsiSXr6GZa9Tq0DMvVSyFrDdK
AH5qHCANOnAcbdv60rbLN2AQcil2MzphwYvMxlLegAOoUYRXP629pCONGlrpYsyt
5fjHVt8XVaUhpm8LRMwnILKaGPwYtthBDVYlXDwS52sRmLpKgrM8e9ijCZ9kj+in
i//2t6veMbdGABuy0sAV3OXabhL4Cc62DzYomBLs3BMf6DMa67jLRw6fuye1Ie8G
L020VQBGyORZUxc2tJN6UNRhty/HwU4w2gTndJnww6TKvj3ob/wQ3m19oPFnegGm
l4zFOucb9fVMA3DLfQdefl4woZSG5iWarrO/DoOJ24jPF87JMqGjLS9EDgdlACqg
MEO5izyukGNlQULz1bdJXbo78Kcto8abKa9ytZRmA/uM0uQRoToaRmVavMBRDANm
84tbQYSp6X9HkMmjzUcpIrutfzYiWH3TMp4Uji97MzJeKMLZE+cyo+4t9C4rf58K
tpGvF75fCn1lujYmZgEnJNdSihL/i/5+qgeAq9Om1KcWLWye+iF50+k2/9yMZbFR
krG84mNeBaMJz+6/OHGW2vSxrlolM7aCwMyr48DhUoBAxs7gqdcdACX/5rDCrdhL
5oTMziZUQ2xDR3CY344mhCqAXi6vqx+5Limn4GX+27Gj0GrjaFsd4jtaeordmKk2
wwqhdjPD1/bXBGCEy09+hi50hCvgDHTmtRlcfGZu5qRJRcnMvJVAJx8xprhOB2Bt
9eZtlZXq7BKrnncHvYhRNl8LehYzVSjFf+89x+1g+I2yqfGD6365aGYYmmX5+qKw
y9tR3nAoRUFwAm/qWP7k3x8vB1Y+AOL0EoWH0/Q0/Uu4nW3YacFvEiI1RUS3d+1o
fmX7cRW8jB6cTMMuhJRbVXg8cxXBSOVLvaGJvPzFeHkEHaAmd+4tGV+LbbzT1Std
w4YuRrtGky/h2SpwjkwJX/8JB5XD0RFb0S4QDPvV6PzVQX6tqWd2g4QhsvDq0VJF
oPZykNGJK35HtF298MYDYbJD/aP0WLo9OFQgbpSwUowolqXodciJx81ZVf1CT8HY
9P6kyOvi5x5l6lf0PkX3gPk/UOc8P+Ab/RL+8Atpj+ygz/z6ZMNnKu0kJ8A6nblD
FE1P5u8ABw2fqocJDP5JVdSpkgKeUI0MIGsEwfETEuYugVlwNhB0fuNcUGzN7Xdp
u3PPYeYY0aGZXQDsr2SszU4wPHuA+9VtHUztdCoL6O0nR4rBPmUUU/sFPGVSMKxg
hIEstW+7xuhlE6YyJxNuzGQUFqRjhGbuwNg8xxehnN6vTw/Y05yOgbYfPt7lEzn/
uFHkI9bRKs+3JlKn+eTS5DW6fJHkqT2b8W6DN1Jrx3spIwad36QG7hoC0Ldbu5I6
PaXinbOtBcOFZ99YCRjNF2p284d51A+W5GWzc4KqwD2ayVblrTydj2aaVXchHJuS
cd4ew7BQnyYyE+pGCWJu9b0y4gAhxY5EedFQTbL6KN2ZBQg7uD67V+glwzwhGZmj
gJVRmE0IdboBA+hLAy48VSefprPCvaNiPyQ7JlAkDXbtT0ZSQ2r1ZcDOnO6xRwRJ
FDPN49QqMfLpQK8X1wCP6cwdcAKQcu3Hoxr+mEgicz/XBdWp1hK+E85uVMfTn8K6
o/7A30B9jpeyKijdlFW+8RH3u3bZh6/cDovrx1W4KoLb93AvurBM3c1JINAwEv+u
1q2iEooQyHC+UIWJKszoe2bVr23kweh1H033fM/o6dwaoMz3C0zK0LiA2aZgXo8e
ZG1Tl6d6tOGeHeTuUXb6ayqLw5CpU8LrqiglNLa+ZuNhLS+IhQWy0NPJ7Xekdsho
pOmyDho6yZwgPiIrxnfC2ykTLGWIwQ0bysQgVEcNwVV6qB4OPdjmJpOR0TZtStBt
OUmgV/pRnWHlQo9tWUhXkNDlAIf80Xei8lR7lKHuKbF0qT7nANUBqwS2B+8v98Lj
xxU1ni8hEhs1YkPg3ObdpYubB2Q72B9C4rOTMGFXOyNL4NeoaadIDZ4+Ru8/EMic
06MqMmHaPXvfXLmxGp5PYsDYdpQ1cERzwp4xJgNcNM870OuPgiR/8Rnlhr/YcHCg
7d6N5MqEIkcrdO5kzHCInYsDSR8NQgqdBTetSbTQoo4hYU/5XnbL4j5i0oPJYY5y
mDs2lm1njzSVesyV2UuTRVbbVy2WpLNMUp0sE/d6edi6qyiRGSCgOVhfDYBm3eh2
SX5SzWC6CnGRZDiYEZvKcfV/ZSqbPZShX6xomLgtL5Q9xQoZFBPx2zA3m+rcdoP4
/m+RCg6oB0/QvilaADpdTDYAlW9W4gatkAcf9yw7urijjGzoumw7RchuTC/2k7BY
EjK5/AEzVdwU2xKToUOGwRdZ0AUcz5PQV3/45GAcEKXyMWT+RNqt9fonfWk0OOsI
iMVf1UfmFwkHqBbftrQcKFxauqbC66YJTkaX1qjvKr1oyDhxBJNHZ+tMo5ahFkxS
cFKKjI762GqJ5+usIyBWV5jgHd4lfmGPx/kZkiXh1uIziTR8ehxlGkiD0Hi2U+yj
E0BgSaWq9BAUUQb1IgHbVIqn6J+9FtQD0Fvzoe8ACW+tRjPm/Yn9rRbyL/jZkY3g
e0gqPLGJa7TTGQYHwQ7Knd9DWoWUeBEf6pcIofTplVSp8HHU4mDzFNMUaFxgrCtk
B9aPYyQ1/ByDpJtJHs3ooH5+/REVTkjI5b4S4X94ekuJZ4HU4O/HDCHOF6QYaPAb
w2zRkIvucWz9QfmLqZX7EybJ4OyLJGMdOIbXoKBMeSzFSO7xhXYE5dVX0fjzhBH+
XIOkprLq1N0DrIEcbkva1iYNl3fTWg6w1DwQ4mUrdng7K1+BO7MVq7Bg7jlsMWoj
jNcwVa0dJG4Se3JIjaay8NlaeDba8y1TWjjXE/GzOz720PcKAd33n3B16nOsixRG
1zrDyWYJSII61Vq3ygIwvQknSySJyjCsHI4YY3gml90nVE0ruPseywy1rxyiZ2JG
sZptfRlFf/H1hiKrOX9NNCjdHp3axdyGQ0d8MwNZv2CksVXWOJZTB5GP++k4F+kl
PHEk7AMyieYu1fbTzq/7Q8S62oQlu55vmnZZaDgyUWHilHBfnQYK9T3sGSuvM/dl
2Jtp87apKk74vH21hyAD14b6AqCzOJfvjrgv+BK9ze/DE+z4WjQVksDZcJHAoY+z
szOwX7F4Hv+V4mvGo3ERRbWy6DZjryP18cr/+p+/dzseVp94FQekJEhmBPcT7SdJ
65u3RwSqlXK7knQW6MLGApNoDhwwO/H8zzAZLdxAQBs4EZ1mV2loijvbj13TcxUC
Kyu3RzJ8WqA+57S+yPD5pqZtPeAGdk7Jbi6ApES/5wBr/QdxCsCAWld3kAFukhWT
zcBeUC7Wyf4k2JuaMeozOp8ePEp+kM1pZ04cnz0sEWT/biqarBnNSwK8H8Q5zecX
c9X/EDfaoOl5YR2YMjUr4CuVDOo5F5twLTaq94B+mWDfCHEaRpkqEK/v45QgDrwh
cfDnbrYrYyYpNALE+ikGao32SpKqCagD8USyAay6CtHvrQt6EaVW0aanekUVUJUW
C/msTXQ7Wl7WuuzQgev+ro7aAukdzMQVNOZiRHbpVoJHqbCZ4jz/dp5bZgvy7Ot4
DrCAZfe/VzDkqALfNYW3bhtWPlPHnxZ2WLq9z5wVZIn5ty65sBX73irnhHCCUXUo
85COUXvIJ2vtT7ahSGKsdy66X8XpxE4pVS6sQ5lqYwr74uylzJZM/pBX4qKz/Xnt
Cmi0TusZp+AGRf3uAtm/TJZQWriQsJgbIV60TSBpYifgDLQv2x5qiWijP7f21TTL
aeqpiaFm5MOMaAE9WRDu0qzc4bfmZkCCyrfE+AttYR4YZj4Vaz5L4cy1VJEw7HPp
vaBO8zC0XJbkatE5gm1pxlnNNV2jo6I334QY62FWpOJ0NE1jWZEoDh5cGgJlvItT
CiNs9gsaDY7Wnlv9GUnw3ZRVQWpalm+sJb9l1/KoHBRY7ucNWNTutQV0Zfyzljzd
iDoPwCesLDyYa8+Nmo6VyGWAGcEQDTn55wR5asMWHGyTpfUjyuyvSkGvTc2ryaES
OUhCu5YohqJ5fJOfuU1eptp45NzZ28LXdTSweqG98mVFdgrM5PH5+RIrdxyv4ORt
MijZ9zV28Ji1OUtNIBYPrzq0qCq0w/fnSf/s2mjUIkI0ssrtX5g01eYAZ4Gg1Wjm
8W5Ua/o9T5i6ClNWaNeUSh54oGPA/GW4F2Bk/iKq979WN6dO4MYE+qvxb89PD6a8
+lHkEwSblFdAcVTyM3bfNIsYOmT4JnFFHltXe+f9uGpt5KTpnc4NdotTGnZvMRfo
yXGjgsMO31E6Ti2b0pde40c8dqiEhk3WYLXiwAhhZRpmFs1JgF28Mb7c/6yMKv/w
+deu/EUHPzlZgdxH/Fl3aj7Frh2pyUJrcTd1Q31YFmpc6AM18ewy1bxgCoiUeUxL
9m/WmBWyk123CRmmMCP+KLsJxLEJl8zMLF+CKxjImH506qUNHv53uaOxCUWAdfcG
JJE8er03hLUXM0+eTisL2aX4RHxx5rq/dcNQ+fLiIgBeie7tfRk4vaDBVLVe0iUO
h8V9qGDOd0Kck7i0BzuoNPCz32yjamOsLtHP9irXso7fEfM5vvaQ+3DkIGaiJuWu
fpjq49lbxrJfmYg9nH5yEN5IJOJrUGiVWAbi1rGj5jXHdHlLAuhyi+eSNcCosCHw
eOIeDznRqEjBt3dcCnzq6VNgWi+FYFJkwujlI/SRgX/LN6PGUG6n4G2kf/Ak1oiE
/UFeKHct6WcK3LhSXGNVheDB65yN9XoOe0V222d5L2jnYciGF0p69dLAyxHCSoeM
Put4Bl1TiX+JvAgQ5FTa/Lw6MzVslvp8+J/5BXVfo+7xSlGKU7cckkcJ8pOj7qeJ
0WfI+31HJWZ4FuL2c9xSf+wQ5xPnZgs8skwNukjiJQKqYbPKfjAv5jaN0lEY3NKV
mD/gBNXht38Qd1VNQZgqVUO+tQ0TRfkh4VeR+vY1xQl7O7TEkRtUiyd2NqGEXFPM
q5O8+VfIpe14wrPSmlp8ORszeFE+OBAjQzYyM3iUx511wgKG0+yfRpn3j6LTAWPY
EeV1FMq/+bW+sKkwrCEs5Ok5FvCqValAF9uiszmiX1QRHBlCExdWmP9TmgrWj1uw
w3DvhOO60gK6QVTWIFzVLTxEbdEffwsIy9j9qn5UepTUP2zgoMyHAw851myJAYUj
7Z1SO2N4ISJy6lFEYOtv3oTR3WgBxxeNAf949a/6vucdCOrcfbhbX2zfDJJ62EHy
H4TN7jyd9sYu0bHoGUfd0LNcvaFGPEY6yO9Ud5eUZSsg2yXE29/z5NrBdavowuxa
EKWNouHU4Z+ZNQiorYzrKfI3XftC+rZkCGEjKspm7EyjdC/AtK9fQLZvUcYkgADg
QUNiKTeGRyxTroiUxVmDSdC26bLoan470GSTPioX7UT+a7RJWOrQqPE1Su9cGV31
ZpdjPjK+ZDdH0ENtuK18DE8Nu+j/JyNUEGOX+NUFPBp5V8DAb6R5UgoK8y3FoGoS
3PqxtehN31aZ4ZDbVfV05Du/y3xFL1IfJJ+Pv0qzSzaFsaZ0EDyMNG2F6+OO/NVL
0JFpsCqTJUupW0FYT/De/9e8T6u7Kh4aSAaLm0fGAEF12qEma1MmeMmHgY63nkgF
YnEkeWmsYLqMxRH/D1P1x6BT8eRzaG6rtu/NojTeNao0ywcGR+aWygXfEglCot78
lxlJ3fQOWYCjl5lMzMBYfikgnwJ1MavFvlZp2jpevCVpmrtrTcsP4C0dCvVhYpac
hLVqkkDmTCB5kJR09jWXie3ImsnYEolplMndvFDr0msdXsq5uE2224ywcDn1MgE4
21nHyk0P1+s4UhVUKfepG6yF5Bj5MAWA+JhKrvHLE/9EeOGaXqr4sYe/zVBgDQMN
V9Sbo+fQR/feT450MY2TNTfafEwbq6xZvvdqqfqQLPoKMBPfAlkqULgJxEnlRgPF
gx9ArIllkdHaByrLdIWMMwzNF7VBrdEUnJRMKhQx2LfM7G2VaNzkeS2rkt2Cn8Ug
6N1GO3RWoT9cW8Os/5ppnnTYKfNF555q0qyUDdIl6X/ltZNVK9WuCGO6Hvw5Bd5A
QtGcC41SPbOPwbFnYytPBhdNrSopxW0G32awryQN/LILtq6w7e8+Fbp0A2DJlBN/
EGGK4XlGaIZT3O5sN254Xk3PFkVK7B04iTk6NYKTOHiQF82d5CE5G68yRdWeGZh9
QxQiBV7ZOpuJpoewE5WjeDkBc0+SYNHBdhpzEbmaMXu8BkRtdsWBHZ5X45XNrb51
7ANqkco+COKsxs0YMisO1q2vhubgTNRoJ2dz2Dkv4pkyKRJKW2krhW4l6gW15fDl
Qd3e/WkMJyuTcikJzWN3C4gWgELi70SsaFKSAJhaeDQRkMnYY51H8nDQ4t+vMIbr
jj4iTJPV43KMQem7KYLKOGmfenRIK+Quj2sn4ozgLOQOcFb87VU/jxm+K6VHS9Le
S48WcYbzkX4TmmXYkJzpMh7HvacQKBW4ImgWgTou+XYX1jF4F7DLXP1yYRNv9OiC
cfEcIR6BTstmS+aNAjZq55tfkvRCGteSn9QhdvDQe9GJuJEVahE3KiHJ9lRfJWiZ
c+iLITiIay9lceAkFQrTZP7q31X1JaDxE+txYKYBDi+3DWrPuUXjd/cosl3NhulS
rfBtyjzDxQi5UeMRmnfnEz7GqCIVHcaLxq4oCr6rGwg8Ryt3u7sY7cn8rWFtGYjs
8r0uYs0MQrkRHJ1vFr1EAg5Vppa/a1rDT3eR8s2yMVINSSV5VvQqi4RH99ljAxBA
xlRSIg/3u1I0baeq0NoT0v9kuuuKqWsdVFVUGOxjgzfZwzgoe5l4cwXyvyAr9UQE
O/4Kb+4MWhKqG6BoxPm26MdIWBd9mTeodWkb1LZtcnAHnH+VsG4XbPbkBsDy5q0U
sZal1pQjmagPp91womprZ4e1wZ/+mUbkKrs1rapW3nto50oLuI+0Rmgk0Gu4bsWa
KZy8WV+5wzR+39mFvY5caYXW1kldJ596sdCsOJUiRxGyJ46Xc8r8FMnWq6J0nKx9
et8wENcHDfTMolv02mGerkL8ozJgYoFiNjbSyb5H51hokYa9oGbPqJHeh0XU9xTt
kiebjXCVntT5Guuy0NuU5U//NWKokLYpS9UXrCLo7bkgBJsgJ8h9+8+EjbRPIqPH
kLKhMSGk+EVLPWWASY5uoWKdcD9vp7E+tJ6Y6rAv5Li5JtyP4d93TIUTmPwt4Vd3
B97YIRWky+xr0MvmLgIQ4Z+4x1J1uBbhWbivMrEzISPoNTx4i4ty1KR4WzSISBk+
TpUg2dkkmIlOysvzLYaRwXDVkYENDOioMuGjkuLf51RSbPbgJ1QLE1YuFOBjL2e0
DP6GFpucs1PPTpVDwzvMWpHgtty1dNegKp8EO0Y8FTd4RMUrLakY1RYY1RTgN2zs
RNzRHPDQh6lQAe+XSkp95qDyNIWld0HP10X6e8qHUPF+5bT4y0QdzUSVgMxLYKnS
i2F5JaumxgCmeRknw4ojBIqRwaGRxgaSmexaObUoMevdCSpnTqAALOSymH2MWHmD
+QoZuHZ9cPi81q2Ex9IzLwuOWH74s7EPqXD/XXK8rDO8N2DcHFgyAePnFkmnwtnC
KrSg0gpg5kixvRCRChZa+ILK5scybJ5kux4IDeDOuCxSEiJocoU8mmM5WtXaRZWZ
gdCYe2H2hIWQasa8roT7cjMbBixJxZloLOJwm1O1AY1X/2dTqr/1yojzAIoNVDFM
HMDbRUJq2oky3AmNxt+NFvhY97FkW3uIoLIQUEyCX9lKTb3foh217nRyVrc475xD
tic8fFXYh/aUd1GAN202RdSbwnUfY+b+aSUFLxm+61DPQf8gv7uIpK147Yesl9jl
QmdAnQ36+oIL7g/rLH0BjgnWXWKeW4vMWKaiGgTWJ/Q4VSwjrq2jyrM+lSPxpVKl
b0gUoBGqwc35Juf8nPIC3jJLqNQFyCxlEKAem4lNXVtOqeoyyW+otFgQ6GMQA+dl
oGbt9LMMDtkmIxxYMsntqYon8+8+IvmNuHG3cRUCZ8ycVHWN4j53cUR5YjnK8+FK
gndKR6zjEsVfl4hfLjRbV9ynRkTJovTD38VB1bxgXzTQRAAhZnlHhE1akWIzs/NR
Kb7BBpZPhRDDErjz8U8kvEK7/IS2D8ZHl+O1zwCS7GGBtm3kLDCywGjocFZPCimS
GtFsMGYsaECIKOCGT71lRabIVOFujsEmJfEmaWKYlQ478hr5AGDpYafYooogyNZr
rhMifqiHQPSSm/DFaKTvQM1fSF0h1CBWlYPTftxF8/2L2FJF1hKG5kbCQq06SsbG
lubgo//ETCbkbzPIiu1ue5i74Zl1k40/E0u6xvnLooD6plJvMo9sYZnwCc8BFKd+
ZUVBTG4m+y8I/3d9T3HqfD0lXeHgRUJP1lwJkJoHpmhTgJLWc+c8uiOdXkStXZRG
CpqmjNVtVudX7i67OO4cTc2+OhQg6H56UkegdhWLmp4li4frx1tqbt2m+LCGvTqs
HYHAmkhnOlp5z67lvT0cpbEgPmvTSghP6LZt7V8dMdqtdZ7yQ7tjPCGTbCfrZsMR
B34As+FJQSXHuWL7y5lVUS9k6YhpPifh3iGrBd6st0LVp2AmnEiT/LZky30RdM/a
9fy21o+gyQmdx+ztDHEyFTTlx0WIQDBXHJoSXyNLmBjB2z+duIj5B+Aps36jGoz0
L2KCgR7Na8/NV/tfs7SU9L42nZuS3/lcAW5vfuVYaVFbS3K8RGjEW5ZxAGZIzGuE
+8jweZ4BiWdu5wIRYif4I0tFvTYhTtFs4MzPfVhrIOFbayQtCcwJoEd2XpU7W31k
PubhCLMqxZ3o7YDNlRvUWNifhFiTYVLttayhd0xG7LP/tu9Ikz/E33J0AmiY6Wle
hut1v9AcNQG5aUWy050iARDt+G5WuUVwUS/2XM+PYpzjIy5bQB5o9NDQ6hjEFfh6
5cIuvyMfmAynMOGamJ3TpE+OVfxhgI/J+xTkPlbXw2PbI4VjKrUKyxfxu8LawHsR
51br11JsfDQrpdMS55BweDDYH33M+S7/FtMPOp4N1UeKiqTdsJaQj0EWlpAbjEi5
wvOkdDtT1lBYqE12C428pM81m7BKJgFTT18b5+9w04PkTZeNTrBPWowAW/yUOJv+
Tyk/oOPgPuzk3B8gNgSjJtK9gADRJBrYy77nSH/r9k71iAh0ltOmpkOBvCpsHYYZ
OBFZHWRoEHcuJ9TelozRCRmauM57YpQdtZV6kOmfk4xasVUuaohVTjb0wYbK5Ixn
ipgZ2vncL2B5Zp8gWlTEspyv6mG+MtBZfcpabbQlphXsz8E01mSgQ3E2WwcdwoDY
dXLisdGXkEn4Tn9uCc/4Q89wS1zcOMoaNpqCGVha5dBZSVuO5ie8Dxh5yPdevPbl
h6RukbVcyBeLuvWe7YUIaloF3fgqiSChSmtn2EkXoNiEiavSY1L0Ytirqjo8V35d
rdOdkWcbSFM1lz7TP3AhVeXnW0qPHGGFdfQOuB7f0bhGUjVwa0Z2aARc1hvDKDaP
MrShy/KXNVMchIPhc5sTlNfgvW4C0qmWwTzPYfrM3tBEvNG02al6m5fIaqgCqYUu
QQkrqPHuGg6xkWD7g7Lwpw1mggEuBeaqMkaGKP8aeDLV8zIFNPikAz3YZ3mUWgbw
/7Qe+QmNniYS+EozsxvXkfSX+ow31QbQStaOcJ/1MAdYf9tYB975Ipw0ARgj2UOL
9F2E/g+BM8paymVx6Nz4FGseLn0vjsfiFw7jeTom5BWhXlAts4EldaZ8CeWy0mMy
ADZlQ5rQGviojdpQl/y+brW8JuxR/EgZ3kMISkoKxwL1QvXT3ITuG81bHkiY/rbr
j8pns51OIWhpn+ted1yMc3C59qMrSq3aoohojWm4yo8KfVkvnjeNPswQFX004v/u
dop6QSUySXyCUHMwbRBGI6IabgTOPiVSabePvWsBtmw1uARzgTtB5O9xEPduUbRg
jLD8BnR0KVzHyKX8D0OEiyR52cbNhBJ9MHEo7d7Ca8UCK+SvckJ6xGQIYYGBA+Zu
ZfkblUoeH6/D+Fon3XZUXfX/AaGBVpV5w8hDv0/WLbZFxe5bW310RwRSrC2LukWy
xtjdwcAvj+8aHk8pFnG26Qn/vidi/KGTxEyHs9MwlfvydyA7U+06Fh8yrTeR+LrX
c4bRJp7fQhIxcBSi6QJjOETFvaHsvm2vz6IOk/80bVCD0r2Qjz8awH712aAYoRIR
KMLXXJ8EMZ/8jRTXyOC3hGGc78GGXpElojr98JLirXJIZWDbGg0TKJN+iBla6Ket
QR/GR0dAjiDV9XeoheZrCfP4AqDGNmIocgPqdb9KlXkSddgsbI2sitytIg5a64hi
9N7PTC1zuoVjMlfVxlodvzPyEWP1217MVUKrgcdJkIXRi2PiA1/IfC/wtNn+2sqZ
wHbixp+TnrEv5jGiizWb4x1xvnbBIU6pJ7ITpTW0IqGEFCy5JdXSpTS6G0srAbkU
BwVnrnbEC/pqAK0jPlaoxsP8C0ZLAZVf6L8CfTCcx4vmpGup3u/Cl0FNWPCFfv3f
fWptw/RBs5lBNvX83zMEj2N9lNaYUcCuQ7XKT1d5Alx+FxGAmZERdiRdro68kFXI
pHMrpCZLvtS5k5EtXnX2I9I6Hsy4TxzpRXeKyauSHz1w6qtC/r0FM8v33kxPfmOy
nSmhXQEYdsS71X/wlv9wrFbyXTNYcQNLQEbi+xGl98O5hklPpT1Dk89fkYvf8m4K
9R/VMJWjbNseQAtV67N5ChEbrUgVCi5Wdi8DOGR2HXmcwxyXuJ2o+/dQoe+gxCHv
g7hh8a8LVVs1IF8oO3BSfKMhz+cyDzYQkaGpYsf7Cf4e9s7xCQYTNlexve5ePG30
l15AgDcF1Lb+DEA/6Qny/TAQ7Exm2CcloCE5MFVeDkGcFoOswNhbZpUfoTnIWpwj
Tzg70EiZ3GDFmXnAtEF9QkfLCQ2KAkPb6Atxjb2/8qN2c5J6SSTeg3jIZOgRPq2p
5bmhOW2eFqatZq3PKUHwLkQ101lB8Ru9MZ3WRPwGcNK0SkGN+FAUb28vu5HTdcar
ZldiCnH1mdbY30LlMVHhKkhn4wJ/+xVtiArnsBj5W7DEdxOIc8KBDVXFwQnjw3eH
DFHlnL6+cDipNCf7L6OXbiEbMdYSp9Kf5sLpd4bsBpI+a8Naw4ZQIXyDgObni/N4
50zmzj6jWGR2A7ufi4ySTs1A7Yr5+JPLI+WsXCv+cYcjo1blHRYEifvltmMrbZ7P
z/02hPZ8a0c80MS6exQ8tpG1eY613Qze/zubdfWsH0CNszBnjegG7NN6sNUlGzZv
s+J96jvnDdW1UFhGmqy4H7HrpS7j1mP7ddVKdFnBv7R4hN/GtjbpWmaMqxW73PwT
082nGpNSK/L+slPI4kdYz1xl9ZCMHjUvdlZWra+iehdTmL1PX98TqtxAVEu0CXdP
kLZwWDXVJfnWlYAx7ZWSQ+ADD8A9z8Qklbc88zNF4OP4ZxErcwPCb6fb0WJE1PqP
DopGg95tuB8V8o0sfJnEb3CUFaaHFnTFp+6a4ZI5zr1wdIunCgCia5lFBR5lF44U
MS5jz3j/o21gJs1ZkgQWeXpunf3SqsYnd6AnyA7YxnPBneTr++M7hbvbXGto+1cY
yRdLTtDh59RrWgprzrofk86sa7uJOJSZal9+0a2QdqSKPjXaFhrmIa4t8b95rz6l
caACGJ9itGVnE2/z5lRTQZLStIVaesUHYdEcJE5V+UwkirrRwYbzfAUzws0HzXSN
5x8hmPnx8jNYeJplmW6tchrT88F4qEEj7EmOTYw38UPmdhk+pkQJzqgy2CxGCUWz
Ll/F2TAR0+ZpwwaXeeQpq1pYbzlSlzPGI05V3FS+frsWKi0gGYY8hGRcPVfzHacP
ewwG78GbDLWMfwHQ8hzF3/OXPzEFxMD0K3EvC8yQjzL2cqOci0mpInFzzPeRzG5/
oMehWX5ZsysRV1I4Bd+CcVeB2MVtueABQswLxdY71zTHwRRSY9MTCdO7/WuLmD7f
LNx2h5yKAFcPYtL/KnfhSbifzYNs8Zfp2YCS8wmiUce3UziSFtAY0NBTEiUvNHEh
8HjHctuQ9wSdmqKbgI59EjtsNgDIjZ22oG2i8bnKTwUiOyvvJ1+XHoPwtDud0z7b
2l3yAFmffYBqI92IsLV/q9+B4mfe8y87yH3fHenCg3or+VeeMJvaFywzExbsE4iQ
Y7lmPDmeDQFQSO99TqkDL4HtzZR4i64G+wF6ArvnzvLvqsA8moHizp3f76BkAV1q
kS7zsLbnjDLLXgdlmSKeX5k9VWj9532AKxie4vZ+B6inSUA+cXv5pRyCBhFLULyx
3iXxNKRfUZTJL+at/6icNWipyqp0N3xv3ort8EYuXBcUqgmQwjp9RIKUvUYTxktl
1l+pYAr/xCMn9QTeJz2+FX/62JSQLvzcMpRTZyI9cNJ7CgcQErM4YFpc7tP0p2ew
7PkM3LK+NmGhAB9obIc5og6clQLfY8gDllRJN7dGfRpcK3CGSjr0qAVVN6tYsw84
XoiYgZS8MfXJjAvYAHfNtDlR1LYGkhqr6/la7fz6PNtAHDG1+VCf2h0lx0uKtSip
awNI+VzoXZLTmUvZUaCb89Om6mjIeclmVBk7qzwYTfnzubCHRgIMmbS7YZc8WX3a
5RhY3sEwmP7ymYUA9+xBeUaPWKvd/m0HD0HsMZ5E4xxTYEOjGneeHxDU8NlBRwnb
82PAVrcqNENORkQxto5YTMyXdwM6LCrFDDA4OH2qSVRA37GgiWfu2kHev3E/EF/5
OQBL/nN9LqqeR0wgJ3kJkS8GRhichy9aIBaKCryGjOqCrXzmVgtjQ9X33CY1puc9
rxU2kbdF4YQxh6t58EepKZEiVeGvKmmDwGHUywnmgjUExE1HS9kghsM9NU/0Xo0/
161Xo+p0M9faket7jtu8TgMGGRoyMkG825z5H+TbSTu+bNBO13jpW1kG81UbMKx0
j1yee2vowQRvaMvrLxo+gevNEh96tS1qxXftaHoBFMCBpQgCf5gWKKOKYJQuuY2T
atwVCO4Y2pH9IHMoCl/ku83OtgRIkmLO67O5dczsJbhKr43j0QKATcRdKpZ2NycD
AfIS7jOd/oic72AV3FSl37Q3hIQYw6/OD2XEucllfSJyIszfjUgpmlJfA0o3KAHl
rQhP2YKUlERJHKW14/cne7oTP/ICYoT6EyAK6m0BLMhB3EStsUbuyk9sZbSjNnzg
lRhiIuE5+ymYu1gJYLwQxyNJoguC91c5HdmYzdfF/GOX+FJZKRFfMKzVeqiRHK+f
3qByxCD5enAHJx9JIFnBSHMEzGQVf6gkP21BIG5ySubt+SocfvNBehW+HZGGrADc
HcOvp38GHi+SltyvNGcCgE8/qGnQc2enSZho1MSj0WUM9a+f0dhaFE4yyKGApl/Z
Pq82p6dVX16SLWB1zBeFZojD6qwNPMI0qQIcBMp4yF2B4bbwZvm8yObHBEKMN8NV
j2Q+pFuER2IzlQ84W4t57zJ1omFrvX/AXIgP3n51sJoeRwzde6JbjaE+/xonOInk
oMTd124co6+/HyJ9NsbGS/LYKK54/vMBj/N3dUKgyNJF/JtCtAippPLXMdV79t4c
pkvkb2f1tjNg94UA8WVc9DGvDrswNOKWgwul+nNQYuOP+nvzD4+l/1nnKT46PJOI
jzsCMwmP6Rjx5ngpYsYhO/huy+cclV3m1uF6GOOhyJFi6+T9IjfYCq1DrQiicGs/
7Vt5sR42d8bUsG2X88hyg4Z4s0/2+92ruZz42gSvxWdm6F/CHMcwNerrvu/nt0wx
z4IZD1MS/bEIwQcBtKiwoslY3VSgxIAV9DhHAwBISGdYf5CDDAVDACKtEyT9j5uk
yALrAFMuBGf0OPpwW1ryU2TH+0RBum+FgC38YbS4dm0P1cUM+HkgDWV7Eb91UlO6
67yqzFJCpaR6SDeH8AKWzeQlzVnCsiKWp8Zlyn0fQm7rRqky/XffGh2OqMX8Ydoz
qSvr9fY8OPheAkZJ+acfWaTmHbZ0iVjNxk0UDqar9t749+9sHsh+qtcyGxYLV26U
KbVTNMuFjNSEgtXYVzVNJ+lxi1orafR7q0QiU4pgQL5v6TcwL+Ihn3+ssR7tjK0u
aFMDvZEn4txWt97nF36qACkcRFdI8jz/5+gwalz3YO9NzULZQ+egXaBtlOSMbcmZ
F/4R6aA8Ecf/mMboDvPXs6ZB8fL06pSIVzGZbyBTHB6ZvMY0iJuIrDLCX4fWJNXD
T92UWSvM6Pe4FV30DIAKSz21kDBo/iXxxnRLgnE6b84rMNqM4KZQH9L3awFSBBuo
+SkX0VTT/GP+Ur3hGPMrhzOnflmTpxBm+4XcLsAyjA9UVXZW3/7w1t/edXOEoGi/
JZOimR81spEfYDhPCjAweSX6CJbddS2JtjYN+E7TfeU8ucFrPch9GRMFZ5sLYh5H
O/uL6aem8orjoPU/OM08mvsafmJUW84zysCGmUu6PANujEz7ghg62x/O+jHsDzOX
a/I1LSUlQd5np80U2p0vEdJT47QpCPLPNFTdsuQbEFJrAIZ6bZfrY30bNQUh3d56
pDoVmRXyHGfsFWyT6mi5X+QM30CEP0Y5tUFKGCDY2UG8Fx4Bg0eUZtea8/GLGoiJ
4HZHcyfHJ2ktqFUHXo+j7w5m9fqG4iPkd/8UUrSxQmLYTDiZY0HdgmSVYWtv5y5b
pwpjLcxZR5JnHQz1IHDMarFY44U+gTfDci4RgZaHkpxu/JvdLsVGJg6f7Gn16agw
X37Dz0gayqLc6P5h9sMKBqnnKBBQ0ZVGXoJfDt2gSFgO26NFZrQLMHz3qoFCYTO1
KSPUdllT7YPgroqq5ajezJjnDVJ4UV7otwM+3XRjtdTMLXJ7vHKZl+vble4BPMkz
OiNCjuKeI9+mtAH9BglXx02uOcbT62B8d7Zr7WtQox0y4O1OTH8qFZ4rYIWRXD//
i07kdxMWdU7iXCjD8N8qiHGV4Aesp/wQLdKm7Px8Ij7CozVu9yNocZnPkZAXni0A
ocb2un9iTp40PNRIoWfFHwyTHthDZwN4MkyO+y57fkPr3OwhP04dR4EpN5TrypnS
eSNyVn3JhWewryacspY3w8HHSm/MeR8+ln3P8VS1BUppEOYd5CddK2mdhlPQmMaA
UiIKzbcsj5M1nWAmL75fdf4t6ja+jdi/MqefQWtIBMKFftqP69cq1qX6V8G/M8wA
jmxqt28blLea52syUJg+nH2FI0z1wXgFe6LoHt9JBoIRKxzFcI2BMqmA3/lvNH3+
sAXSDo/2DWkd/ochn9cz0z7sfzQ2nR/Aps292SATzGj2qtlHM62I5XuMo7MWjW5S
SE7iP/Gmbga4a/Rg1Y8bEQ9rGAi+YWM5oKaXik8R+COj90hG3/l8gWY50OvYmeV6
t6K5alpNVbOwZrs4hys6XDewsPPgQbHA5Vw/hksLZwfqkzepGapWwjD71JrUDmwB
zzWmXR3lksM5VnLL98w8OGaItz92YLG+uTDon7F4YhpGW5CV+L2MhRg5biIK7yGF
btrbn24aEu5IPLJDgJl9YAIT+uJheRq6TdUmqO7Uj8PTgBT+8Zur7hTFibiMVYy8
w2RJEnclU9v56hkHTdLsWgrZmgEhI7JO04F+TOfZVEKhrYUY/E6uozTdJSxrRfcq
/Oz/Csdu78zZcse8oWcnzdlKb7F/OfGATkBjk7EoeKm1tN5JLCORjQ1hw/wW4Cg7
68gSCHFodujm3++9WVr+nBzuok78HdXXIk0NQSgxN9Vxu/DzWOx+X5625MH8E3Wy
Xe6U1RTewo9k8VgBlbPlodlTArvsXZMBRWUyfmJ++uQvvNzOswWk4nbGU47eyhBo
FfxYNsDB46BZBUXrmnKNK/L3sp/uWhFLV9R3vINOm+5+mZkZzLeRtCer5yQ9vUPx
TDL1j9Qu90MHGHO/Cj6ZZCoa7n661lfUev/GRvq976P159J/+ZZ9kWRzNsHfH/El
AKbb0nCQZZNzm3yUXWr4B6Rq0bW02bpP70rtVKNertr4FOqKRBEoXn9eqovFBi+U
NKhkq41QbUgpTn61qu6q7u3QCgKVfpcvuknfSXooaQx53mHA2wZgSTCqYESYUmQF
nCO3iWCPKVai02NHxtbCk0HNuP7RwSf9R7U3EgX1o0gOIRMOrscH13ab+Z5S6PKv
2uzdz2TPVUnDZLQ93/+iFeo1ILWLq0gT0vha0ZWSYzUEFPkkflzolfjAWFL20Voq
5bXofSNZJ3Q3+RU2WXRWuotETviBfK9PLouBLJP7gcEahUxeRgLTwAcayURfaV3U
qL0xZxbcRpN9ZSdx2q/aGYUV0ZSwcPcF3uy7PgLWjeAdNYYnwcL1imk8rk2ZRe3t
2agiiwhiPguulTWNmQE1zvKwEY5X8v2InsMPfuhCxT1wZxAMuR1bxWERDolsu37N
WNXFhRlkSvuNEgSmo6urn6Seapx7lXAih7JVPee5ElQVVV81vRy2nAxJajEPVYjs
aaSGdu1xzdoQOnux2u7oRPQ4W0rZR7k8OyU0vaeHccgAjVkIU1Apt1lyxxvieUFg
taa1jVUQEaQC/UIT/RMcF7AmREXE/RLR4NyB0f1ha8KDkKwwCO3AT42ghUgIEdnD
2Z4pOEuf1XNXOXVuYb8dRqnYBcVg0h1Sj4arcX1/9SKjhVDIpIoHUSC1cpNr+mZw
IEqUCxsYbuxftUkeC3DGvkqZG5qiP+9mHJJ8w/sZd4npLQM6U6iNavfY42/pLpCn
YBA+AbNkiHfJMi81QDgeASfxf/UETzJoYGq44Z8FuiuIf0FYJGtfwTertA8jZPtG
kW5smSCSRBYHMTGkk02GiumkmAf3Vu29z/jZhIokcSNcsEpCAH2xhhgN7QXQeAGW
Pe9odzSfRE6UNE2SOmnnw2L28M69fQ7rXM8OQ2bIE8p1bMTMyDD8ObWTJDPRbfBi
ZVEzt/XIcPIhoAD3vcu4Rkm9qRSNWwRnnNCToLRJWQ4YXgXCCZquwQj4oWfSMSIh
OVQkN92tn3i98QxVY0I/+ZiPt6dL4Dq9ityF+r2OEScGJxnObjd+4smEdoI27xiH
9aUw5fcjffnDjglgV63TuPFxFBSNsOnUGX8jKEjFwNBj/a9Ul2K/uVjhM6Q9Gkev
dwwMGec8Ht6mkLc68kcXRv0EF1VJlHkCuHyJfXAxxKhUOfRPpfQJEn3tR51NbI1s
rwkY7rvpVD+YO/WjEtizc9EVEe6MBL7x24gQL30QiL9Pod7M0yOCaT2LuPmlPXLu
P8LySnx7RnJ7Xij6nZp3a3L9HcA56gykoXh8ZFm0bIU8gWsNK6jcjn5owRnI92zk
J3UCAw0gz8EJEhVAH6DWcsYnAatZDSktzmOzTdSLyNqXLZykpI1H1Eo6gjS8at+/
Cjtx+NDSe9AP9diSezzXlmFh22ysYyogWzw+pEIYEjy6cDgOiplO96YkL5d8qHP+
0ppkmBbooP3mq4+vN9x17dXmjQANOoJOqJekfYOlczGIXZV/a64h9Jxp1PeQAHGv
5Am2oc2oYrFcg681t/g4jR2lR8kwksekLc9j5qUF77LsIRiGlkyEdb2yZW+48T1C
JyaMDhX6VRKkunZoZql0VOWlWfriVV+3LL2+mbCucO52OoTsPB2etx37jnwYQBMe
U33McqhKUDGQ99UwwgL27IA1hcGu9oy2qX1vdxibQhhvLd9pBN31llGCH8cmrLSy
BQrSFRzsV/2eAx85VzYwa47w5BDblwD5q7L1AwMsF/rJthtkWIylOZi4/1vPqKse
0lPn2hraVhAmLNSJGiYYZN9N3qXUW7iO4PIAYrEkPYyLJDpDZPl07bduj+ga4+r5
hpy66UISyl3bUSrha8eaBttqvgKP5KPud9DOcor0wQBJqp4JWB4eP3wjBrI0rtBK
vFBym/KvrmAuhwCvq17yUznFI3AMeIx3FLN27754C3K+vLsKMwYXgMn9EvYHPw41
R4aEOQgidrCNNaAg8At2oJhraG5Puw/HWKZrcAH7J3lAxSu4MDAooApEXuIbWIqo
fvADcrrhI7MbojBf0UCCSOoacFkaIY/lqvIl47e8Zv/6fv1QH0mVmbqMc/8xQvin
sEEV/9wL9nNVT4/Ij8smqwFF5PetyOllZ9llehie34E4JRV0Lhj91EixBaC0YZNk
3HN3pHrdCzusbzVKLjrKac+p9SXNa7d3PmWQ82blG1w/WSKh4d6i+ac46JJ3hphk
PCSa8eriXYKWevSh1SLTRqZKIa4xQnPrJ/3TStSnrlJzSxu55NVzbkTOhxprIC+D
sVWsjkN7sPIddY8ZLysqF8KCOfSDJHk2JEdRDsvf4TOpLrS69Mtj47ehClzx3q5t
M2ToKOSyH9JkopExyQ92BPuWkrFd85PUQfaKoF6J6oths7wbXYaGeSZppgYewhEO
1riMlh/vttKc7x6vUxyUii1P+a930pSSyblu9btgfD0VCFivnOPKwFGZ084y/0k4
TQV96fDB0UdIQnMrjGG5/bVMHUuv9ZnLY7HapzmBjBTSECDO8Zvjjso2I7lAlzcx
Tr9J6jKPGiixR2Od/GoT2SFSHhJC+sy5LAvkqfoZg0mdDhi10gqmUhrMqDkzoF39
OzuikSncQocSN+mJE2Ao4LekkFVgGsjnAT6GWKEA4+67LnF2dwgHq5sOpb43u0dE
8TXJ+xP4kENQ6ueGgqeXm+TOIoOUei8VTz1KTdK/Rqkb3tb9zF8RLydYTYn08nEj
Tvf6mKYS7/2kEEFIFZc8g1wLEbqOJCrov9B60KyohNkvf60jTlwpLbNkUSh4aOnS
gO1gd7d4TPfGx998NkfNfcLB3dyXcct3a12Bo1rcqJ15MdlYH0D1tUh9GKiqOcKf
QZiKQxc4IjU1ilJKJeGS6sqY7Fk5MylfwRo6sMwsJvh/LqqZ4r3aQZ+TjO8Yogu0
BTw//iIrVNWEDDUjdb7W1In6t74VgzQfnyKJU3URgIbggTJDU9wOGYuXJ2VhUBG/
8PDyUJf+hmqeL4Hg+ZbM4uJ7flMibjewpx7gEeSqPJzGvciKCUmDaLrmMM1y3/bP
meFCpvfOBHjf1y7tBtzdwUEfBQNG3GZwETfdBF+FVce5GotllWBWOJtwWvrgaLo3
zEQ1flL2Tmrxgrl7ZHutJolb8jcSWw25E3M2FLCV6ilDOPBgvEQK9bTKdujrRvtT
nwk8geOxmLi57P8Punt02f5FwmPcQQ9jbVbQBCaXJe8SSEQR3TpWH+aBVTCnGB+h
JUtHytbTfVUE/h9xMi5I6waWCJWinuDtezhwGGHibz3HwFMsN9AXLMqpR7UAnN64
HhNknraYKGIPj+1pKVq67xZgMXH86r8yYsqPL9GUiLKdoua3cxBu9cD3JmvdMGNy
nnpj0+bTj9YN8IoNwJbo9keY8OuU0eZ3Pos3mH9RGgjvnpG91ZuuVcjC0a7gzk1W
ptEtNTJcvAJXyX7unymSP2SGi4U14zY76CuuKOFssDseFvuy5dVHQ12muN8sDohx
a5sn/Nxld3SN7y+Hp3YA4bLDp1RQq3izRdoDAcFLyLIyUmiZf6ZbWg71MEVoJm6a
x4GV0zo5vXWSn6SrAYMZal6xSymJb2Uz81Ul2x7Y+w2GpYXSGq5SmuDd/EVjng7y
eLZfU1wBahRrR/XaXyH321L/KuFsNC7iCMszaMBMnEgE7GfmC1Ah00PyW7SjIGPQ
2zave38GYjfrrJqkBfwf2cPxy+Jr43BnLZb04esFg8SjvK1dXofVqkWfU/nSL78h
8x2ZYWyP2Q2bwqvaaYTT9KDCfuHnGohmU6vtLyUl58GwfPp1AE2/ZJQNIwC2W7Cx
8EVNof1mq700h0JIsMktQ3IlVV3dxDhoTgyag5J3T0ce3n0N1f1L0zkN+k8AH1nQ
1Yx3zetjk8BqLfwecaU6rwxFHSFODpsdt4qn9zVCk9pe1vE5zyJxThXx9XF/Mg8y
t1h4+9Lxgzo6a+cUQIWRh1uvkMkCIxNw4MTx3VI6yGknwKVXQm1PzH7wXfyD1yj7
o58f/7qi1LFT2wcb+vIOKZEv3YvHLnsg3E0Y7rg+K5XLUKxRh/+Mr+HfY2emRRRf
5bS4iej+ORHEfqGXMI003smAxTtbWuCqxMIptvdUx26gucbYKD0bzA9E0ayWcN6W
nk9ccQC/48RpeRt6+78KMJaWgPLj0KIaUiqR2JBNgoC2+TMbToNs9sUXOmgpQJTt
0RL97h8az5ouPh8i+UOghf6a0r5pKuNP2ecdJOK+0HySJeiv1yH7IbqyM8r7rrkq
tciIWxEY5PI2wbjgAKyyN1vPquPs8vBfEgTgHelMAfAVA4XsiGpU/u3IH0ysQD7b
OXERAdNKwLKDLrfGOhgHsOPSgrcEVBh9EyrWirNimWhrl5SmVEhfSX1eNn/UglcK
oP6FArg7Jje3Ovwc4hJGYQc4LrjpnOUnqYERf7svzdlB3QVqm98QoUQaw9Cay/qg
JSKDDDR7pNKmPN9eo64gmrfyvRw2xqSKYgNfTR/bthCi8OznAMOVHVqisA2fLsgd
Ui57rWvbkCeD/OFem0kV5y2aQlW3XmiGttyfo2kdac8W8FWYumrjB6jMgXAgyGxR
iOBsrw9Pn9cQjN3SwEkU/2+DjRuSbOFeSoimTsuZfoPbBX+PbM/YvwaKSNyXKVKU
+KvttmnlTalbgI3/HcceqrEyqYdT4SVjYc7SBDwwdBpZ/i/I2cBYqkbpQT8tPgcT
JQgYkiJV7P2jgRo5H3kGE4u8Tpm7SxXhNWP75mvCVrYpAlH3UUyILnTCvrbwivfu
t/r8QPpv2t7IbZ3kN5X2+VvlvVr0R9fnrqF2Sm0AqJeECU6k5jTmzkQrR2gx7AMH
or6MPUOETbZOMyyy58ej1+cRDQfjoLw+FBJT414HcJ/vlBfynV1R1lMx2SMipXp0
b0kD7Bl71O/ojZcrN/Vr5Brbs1JTzUiTmeaAHTPUCt6XuKkFcOWDMJdHdQih1P5w
LYpgaCdZlwFoY+uDMk3SsVayqWygnLaOmPlSGeSKJ3qYJARChhJZzyCO9Xhm1wyU
txWsDKKG1qlSUxYNXJTIYV/Vzg4XcEYl9lyPEpxkGMo05DuSYwTXv7b70HrtmN/v
cKi+lenldPWgBD3REarDeLlT5g2/yMEk2lgViPVI02XyB9xIpRY0IsDXOvNMX7L2
+I0S8eNwijujoeQqtb6UodDx0dVO2jS2+5QZ+pUG5Xml9d4SY4utuUPvrRuIjiGG
GMuVpM6OedSYEUUXiNqe++aqWioaYDzExz3JYgx46RiRyr5WgW1Rt8JwmeuF/QCc
UyReVOLEQoqas2M+rtO7G6K6ayB8TQI4L/Cg83lUhhwW5NIDOWJkqmQznFCPyHgM
BW14qgoXMBwo+V11J/w7TDPAOzKeGo7jSaVotCJsspddPPQnm16xEZeDxW0uxBG6
vpkT2WfNw92L3kymRHA4WTLuSq5mFHRS1zZuw6WLry6Z7ns+i2mGvh5TSM0JS+rw
jivTFSOMo18kbQ48wfIKYjJlY7irvOAuYkb3By4DKjA2uxEQNFwdz4Nze77Kbq4g
On23xCi5Ix8egrzFK+zz1oXjjciJT6NfWdTedRdrrPJNGf5W0FJxipSuX3hS8LD5
WrANobKI61W6CQvoIJEQj3iTB6UxA6IKWZ2EknKF3YCC5Flbe/DQWpjU1kTNbPRw
YZZGmNZMr/WRC5oi2YfT96MQ8uFV3I8w75MQ3RNRrTGcl6ehSzqn12tgB8jnqx3A
XwUhp4oQDTxlZXzgNjkha0zqHRu1oPfB19I8S897h6mYXryCae/R/gcTQe/nPwbx
utRhHQCton4DFUmI1ecbwTHTLdZteWCOxP10Z9Rj6Fl6Q7hRar/+GnpDS5jHAvQW
0mCKggBbmM3nai5XTGNA28nvhBs0AiR88ODLtZQbLXLtbAcNZxQx6/TWPe892/8F
V/A7nK7PHauzrDLhafjSoCP3krNs+OVinreNrCwrP+5L3aO18d4c7LaEwBdMStrT
1+nll4LfQZ9Sp4r6Ud0NW8ZbvQaYVcIhtFZTH7leZBsBJQNsHB8n2S8JXWlppAX2
s7xBeJb3iKPgyTqFxviysIg1tr/4Uy5LhEH1aEsV9FUmvfy9ekjhWZVsnn3D+NL9
lIgwUUeT8AMS6vwrq4619cceHni+cm3uaw1x9pJHtPg6LRko4ImmVddIoDC6oLkI
zIy8QFSzhClTvxb9b/FpeXnvJDG98ilWzc0WRJ7GX2GqAY9dQngym5FzS1/FhEag
GomMV6GdPOnRF620C5MnDy3+syxlMemQkpdhpRIvdB5UAkI1GyuuKYPzTDJyzBmZ
7m3PJkmZY3b6TaziJD50cMfUCM4mdCTnW9VW2X/HtlgDuvwhXxp/Rgk2OpdnWdR7
dmWPsn32MdkmXbrf/Osy3vDCghhjl6zB8g01rZxOmqdDe5qMJglAc2+GYP7dcUNn
zJ/QH5hrsyT0/ECKvuMZhAB2b4AcpQARVBRP/4rAovJEf+RRuhZbVDN7xdApc2C+
fqdmjlnWPHnrPd6NckCG53FHlmJ2OReMvPjXl2YPq5GAJWoOGnIs6IYP3+TtpXF0
Ajo99SoYBO7LOspbovtW7sWeJAfOsLPIHt2Rg9GsolbDwXoyp52uLumjqEI/NRfh
/WJ6m0k2Xom6wBHX/3+7bgVtYXOW3ZZZqq2BOtXxq+Y0i2MWtkLPRL468n1oSHFj
5Nzds0YRK7gfRpXkMWg6k7RdxIXOfdNqP960UxcIumP+zXoBX4mu5OTXFgdLaQB+
lzCTP3j2nv3bNKX1Opgg1z3EkmpW5JCOejUARomrilHSd0PaMhYailKIdDehfpKg
5FknFoR+qJZugE1dWJJ2jzFXBieYpzD4uDs8eGUwPVdMkBOH5olb+Hk+se+wFeYn
znLUdUcW2IR0onNvEgtN2dx+srmXFAJizn/vXVaMbOX54dqQtVfMfFQJ+eb2JYtW
JS9tEiDIATt6Z/dp+Zm0FH8igQafgk60lKuK6wGB4VLfPpL30iF4dy2uCJZKWcGv
XBlj2S/+JpCg8XJ+r1FTeJcQHQ/es3neYAaerWluiSQFkak9xEGzp+rhy1KlkxvG
ExxlRrr2ScbPxD7qS279Wv0Dp9/aD4s2DwF/qCQRPGVXvgo0h0VPUf5RHGgFM4z9
47cYCnSZR7yc8JrElb6bq8Q0BqKa7WZHu2RS6iz/EZm3kZM9vMblTq9jcGLApxpq
IvBPLf7SEgdOUtGp70jsjblIESKsrq39WFm9u6nYyoIWH3o28L2FwBnsj46TkjQF
Lz1ibitQD9Z16GBYUs08BTUlkKeDSvUutul4FgyfUR3mIZNZhY3iOabHg5rO+5Wq
PQ2zdUY4dFR8s9DqXosIhPfhcrKYHeNEzDq3sFchRZGOt+kV/vg/ls2dXHF1IsHk
rmZNG3XOeGZNxVxXGqrzacwKow7Y1QWxqMR3QK9JcAAN8q5kLm2JfoNybgWbHEOJ
SAkGXzFbCTnCn4qBykLbHJVxmJg6iVIZrqAg+OC1czjHULKIGeOMEwudAcdjr27C
Xrf+KPaW7AVdyC/nJsEdWDX3RI/4zMLGYygnaobj7C056CqYkX8cKqe+UmkPGN/J
cP/oPdxC+2GXD4aAW3W+6Ql8By+Do97vkhNb9MQmw5mZsuuMIYr7pyjtHDxneU6I
gQow2PhVyzoohsBicMRG9Knwf4LQ0mAoyw1SiF2iupoW1nrxYF2QZtWIIHxcIhch
RSBLa9qlZu8K38w557JEkkmQsals6SDVlDkmjOlxWK2ftlrIZYasvuIFYjEwVdxT
DPA9DuT/XIe1L24jxyhfBAhicPFAQ5v0nUB7D5Z5XE4TiMcBj/wxBfLQQVWts5Ha
staCDFUx15Knn9zdkDPkAKg8ejMlIeiY3UQiWjSNC2D8H8KnkN6Ld+prLUCBofnC
nYkPW+o4EKVFNIkYGmUWwDZeABXdzz9rqzOmnsvUKoPpV26s5jkCyOROcj0vWmSP
SYxM+GS8+uLBh6ev1wG/mqnns48UJKeLwXcOVv03d+pB4lYyHR5qAqGcc47sUXyn
kPbT6Ahrjdt2oRpQt1zdjYhgoZV2cz2hyfQF4R7nQ86IUoe7dUeoVRQ7/QaPg4XS
nrkd+AAQaoTpsgwl5+nuGlEAGW0a854cxjllzXw1gph+G+V93KQq7nevsJB4OjJF
AOzf8FA7Q3iHSBzVZz70VnoB0fab542NJ0RLxfgPov/p9ipcsCE3wjr8ni9Y+JI8
ocs4+1E0niNeeP3iFQcwDTeCyB5NQaQA/ezuCjk1KWmT3md4DFUr1LpFxwai3O0X
4lZidQqKub0CKl3qf2WDQX1CUUkqNKsjOXq8F1jTJtjGIZqRC0N9fx0B5hSryXpe
v/s63JpMp6Z9p7XoaYcFFST/fM3tQbJKF3c5N31RgTL4Nz7Ac3BTeQBEFTmYeNRP
7cXiZlx+734bzLskZ1lK/NNfh+paOBrm0XdHQkhOVhVtXDEasewmnqpOD47QMo//
c2yYGlmtdeF2U6EyuEJkG8jQcE8rFQ1KcYdR2Ex8T7WdpMrjkbZtUhKsHridnfKN
CtZd2maOEETWjNjX/6Hp9af7C5pdQT/6IWexbXvUJJj78E+1Tfws1tY/lTZNcyrW
aD0y39mjz7xX5pp1ZrPf4M8WTacf/FoBUhXUF7lMoCp6HaTF6UKdjf1wCBPDdhop
wvTzJ4SOJJ8M//QNckytso8MftY9tx2itEkeKoCcKms0pJ9w1MpwvGkP4IAY5OzB
gz8a14iDfvSvYwJvhsha5ZLlutfAu5J9YLuCYXFkklbSG5MAqPoDRs7xlxODF/NX
kHZt+8SZ3EeAJrAWYmo5Y83PXpH5o5CYx/8xSD13WfpYGwCK4+wjGWsnqHqxeFA9
8rzHACjemsryl4vy1hlzxPamdLYHXOdxmOnah+r17hRVuEpmPZZTWJsdXGPoD215
lzb00gKhQjSdD+wNxURJEgCd8s6ylJaD4TB7Y3qaN8S8ndRAuycURCz4792c6IOl
GrjCQ0WKkkY+4OtzUIYfmT5iugUVVGUNU3uDWc7Bf2hh2C3UYsWcgzCHpmCKYd48
Jp4Ho5ho0faFZ/XdNavxKGCn6abRNjzIbfyuuNTQHWmqwITs/6IpqxXu9cocuZZW
37O/RyUkzzVazhl56h1f4wNynRvl/kvpdAtjVyM64EwDBPEzq/V5J2vBA72Gs3Hd
qF0wZ81gHCCVw1zTVwt2Ux+S8k166jLD50s4BixseNBTpd9ZJOUENnwj6rpbHktM
BPFIHCZNZ1AC2MH2eBRErqEmwBjWLmLXp8+OgD4ryFesZRU9dxnbRTh5pZ29AX8P
wQRoeFwHCwy9VTz3dVld2SHwuk16flxCympFhYXdHRLhqrdUkl2jJ5qbcdmgi5cl
cuyAZB2yZT6equ+7aV+jSUQwMRHX20D9vcCOi2MPMvzdZBjMXfpofS8SzK3GyoDM
Vzs3JykZAvdgn+mFbW+lxVl6+Sr8I0GN5Kcf5RyZ/bgDL98SaknVCcNN5ftUUQh9
XHGelLf4qRnBxDoifDdehTTmgUA0ZNoVBIA/WWSGWpRZl3yJYWR4mvtwbOhDShgZ
lmYjwbzhiqSHjFqf61GivNmkvnCDgTGAUPlSgJ0QHB08L1fRmaTO/ThNvD3VAOkE
VFfz43rKtJKCHpxUHEQdjGAtRbGdhfgdQapok4jcRmJBCkvC2bgWChAfofssGsgw
TPfK+slfGXGdpXBXgqn11XIuVy8Apdt2jJLMd6XS2kVOhU7dgA/uEWYj1slNCSCW
M5XgGvP8an53kKzJAm4nG5+QWZSwiJ+q8KkqHW37ux/JO/0dx/Y3aOCl5RtnhVbv
eCoqCC8zA+wh4L64SDk0jZaWJUC7o6Tl0PJU9Gi017aj2EgJs4YTRLwl9yDt0Ps7
VA4Zzg/GPy+hFI0z327v7uz4oCcTqEPSjZV/yCTTDmTB8CegkNYMECCn5Jj6pkq3
XawgvYWS7BVIW0lspGuARJZOWS0mkABvbkv+IcDFzK8avHO0zD7x3KP00uoUtoe5
+dE+Tp9dEkKOtNx+LOXGDh8ZEkOMKUg5yvHBeEOmKwzr5jSkQsGSos6ko9eRPJNG
OTt1IWuX0IkblnQ/HusidF0P8GdKaHV6eXju1w1Y57+a4CDBRXcqpNPEGTWIMt/i
OGjidJb1pWkSz4qkYiy7SUljKrY0TQLEL7xVm/kG+Fnpvy6GtENYxTqYRNxYuL+Q
Y30rNQ9G7o/3nZQ5U6vE1CTBh02NSHxepSF/nJasgPshlPk4JQVIlOycMAjSnB2d
0R200Y0SxM/itDhSp21KAd9K5eccsZrZVPv6P+l3zQwacNNwnn4mXp9TKaOqGOUN
EtkqH18hHM2ax2Mc1oBr4V+fmAIf4F05X6fak2gGvVEU0SWCvM3DHR4NrzyZgPF5
cDktpKQPqR5BsPSSrL4UtV67eGK5sDUcHd6UI+yoJf3DuUU7Uc6wK+w4BHMhXghW
gIWCdfE75w1FgctX7p3giRPc0cffaDgOsa/3RuJ0a8FfN81tBEH/mf+M8H4VSSt3
2R3Se2wIxttjca10ko+L8hWdJFmMj8fH9eBcGR2FSQVwNUafLh34MxMmAistUcGV
R2Yf+SABBMdbKBMmI4zeDLlfe7KB6xBO5crA4khr8xzxxkF6+EI+9XlB8o2NXAtL
+Xbf6BC0B5yGMprAXRRf1W+DPSlecobCBT+GgbrM+pXzJuJ4jHQnGr6jHiHNXa9S
58Ca8awdRTwzZuy9skQ04IxxVw2UqLgmvuLw0x3CnGGlK+CiBfiIZpl2RZg275SW
WX6HVn6XdLyGqEU8USjBl3J59EZvuvjqqnBfwJnrGnNT0avX3iZX7/VkN+wyZyc+
cQoVwfNuQMHCYpEZOkiacXWYc+obIzDdn0XmKdkBBXXcrhSvXX14Jv4RRqPr3W7e
z7kYU6+LLGdTx4migcsJFKcFGQ7iC+SbC/l2UknV5B+BNnUc03Hf/GYtrzJWJCgd
Px342pcd+w5Semyx8QSudJ4lH6cOeRjaxVR/c04rm7uYhfnrYgkXTdPq7ybaZRvc
ISz7WfB0j/Mg9YTdGWW6TAiLJ2/SYoKg86SsvMbxkPx1ksumeGcsSw/rdR3Tah5t
YGo78GW0bHlFv+53YEi6NqxFikgWAM6NRVCWUigKrwkZAR8IYnRoomyVZFFsXObX
Ylb74WQKmajWOMUmGnZ/TAs5uEwCppnoxqV5ZAtHqldmePwi2Dsc0hfPZbA5ptpA
3VyWpha3wfvPhy5LsGMuCqCUMpgRZ5pS5iBxnw0JgBPHwLmu5sRySoo5VPamVwlM
+y+Fwk1yKGQT1eta0BsP6zxboQ7OaVYy21+I0SrFKYxARQI7F9Zev6BbMSqtllYq
ldyVu3VgORzOWUMQdWV04IXyUfjOsWNE9V0SIK8GlGbkr6xqNedEx4I8wAmCqckD
/a2ER7orHD8MSZeKHOzk4G1K3+DrBlB/nwf/HQzx9S/qaMoqO6l6KxRO3EtiMNKY
sBoBNid7FmzSE4Y2FFEtnkB1hwfps41SJTuqfI81EdYbPOCj1j7FMblZS8bS3HKB
idr/Oo/oEl099X4rsnkJyqe17ewHb28TdwB3lqkHvQ5Qwjmi3KSeI5MI9KI+aGuQ
J9MNGhlWC7dXeN/4mrKIK9iPIk8K0smwO0kIuPtJAbBMVkZn0cYS8Bp+0+/ZJzw3
jTHxLKgBQ6YXfGNKO2lnkmCzL/oB62OOEg4IZVPLOg99HsuyQANHso1qg/ms2tbx
SEqaSZ8O3KCmKibqFrLNfKqWwCpkpKTfhDT9yccE/n0Awbzm5h6pbFxOvL+M09fg
RRYH6EJfGhSFi8k/VwxUxnRSptB7DemEVN/2oF8m8auLWM3WBfsEabimWDj/URzY
zj4uZxAWmUeios5oka9cguWWN02egoPc4x4F/My7N/DSf8qeokqIEAqmofvKGtcN
9vzRoSd2QTqvSJ8C56dFwPeyjss3KYOpKQmuhg8vtMbiyKp+w6CE01QsbFS6REJt
YktAJSnzGm+oyNaASYlt4FJ1eqiOas+QOHrjP6Y6M4oq7OZ1avL7QSJrL7LrqRKQ
+b1ikAJiwSesuF8mXZWLiytppdLFf3TQMdhi4MLDpx6uEtLNm9N/URi1ZasxTkXP
yfytBxL0kodHuvFGlzOVNEfNVz4uAreA/8xwsw+b8XSUtWzGcdPWmF+kGxmeqT85
9FdeT8ElFqrsTzwwSUhrMREh/2WryUTgeo5NV0/KU3gZGayysHTXuNTcnaAvj3AS
PbqWw7JbgnEhs0faPuHndDC44r6aBstZ5pDf6Tku6J9V7uvj8+4+spX8pxVZirwM
hAh+uu30cN5QNJ9w8yBg6vplvqs3JWHx/y1hf8i+HFcMrLYdY4WgiI7jJOu1BSf5
3RFf9MtAUStaf1waNUeG2/u+C8OUPXg/wcrG8VLvbjqg8tz5dOVWju8l4FdOjWY9
Zronp2x8TORppQs11o+/CEHxJUYDnuhyru0UfKFL0m2fhBY++XN49P2FSqekktOC
mnWTDJ3mPb6wntmJ0rllGyNZBlX7XeyMJdIpQ73RrxRcBTW8k3PCaRsb1FZiNFRN
17eMA2TWuedHPG9BKnSo45vN4n2keDZS1EVueQcr8+J7E11WpkPQSsKGNu1JdNF+
sE9xjHdk7fpm72+lDGMdpDu2TTdtOGFHqX6KsxFJqjZsyiu0FnFucr6MYyFizPcB
T2op+x35A2HmqaAkQAcAKfV94ZkhSUJvEnOs3PeyDuHn/l+aIfqr6U1k3u5ltKuj
UytOR8up9iL5ab/DbRQDTxc0nhA3QiPuN9CAdizQfzQfE41mfPOI9HQZYZoQ8XzD
Vvbm9MF+xyqx+2T1FPsQYvBXS1EHj5M3qc4fFCROEMoM7uVorvy0urBPJ1wnkVOt
T1xjp115PiCSqNoEY4bsFX1nOr+Cbd6WRz8F/r40NpXLycpXTwfdinxT90WF5Jt9
X8PfLt1GTrI3UnVNyalXtSUhXS6YJjdoOV0P1a3mj8ZmKkgR+P9gIL/5UvWBzQ9B
PSovC6X5ks2HarvgluIsuOJZjstI4tEtSaur6JQarqMbjN8LBNnkD5EFu0zDLQuH
XAz4V7lTNnbKhT3RtodFQ93AsmIvfCQq603Wbl9UjH5k8Z6LI1tx8M5RD6uNFapq
iXxM98tDP2beCBqmcn2tGd9kn722DFg/ZATvAuXfxNEANsUmN0Jvxio3iWwZ8yd2
H43tcYXzgcc96eoFxZD84q5rLgB/nqGAReabLW4D0WROSqyenUGYXRf3NsfiAEOD
eB2bhRTvm2s0hE98M06Z7i7QrqnnWmjTCzYyQj1f9ZHSQc+AEkAjiEo3/mlGeijZ
bShkO+i+fxon4sfkM2rdjyNzeAVrrMjp/R1V31jOePCz/mbpB5wOl7qcJQxAIgFl
nYYjmtTpvFFEJJOgLPfgNigrACq5Smu6ElgwNLLilUGq8bGIrf+KgKmLVehzs/xj
c7jjhsuNPwHF2lbyCtDJ5pjMXDDbXG/6I0jAYBw5QeYEVQhl/3tvSLhh+1twJNnx
J2ZkQGzgKUIk2dEOZzxcBwgz7kRI2O4Vj4U5Oyj7d+rTovHC2/7S2DvvvN1O/n/D
tVY0DsTtDvt+u2S+IsatpN7db4hU4n95IWsJ6D3MMaY3fkoTPskb5CFDGydDX8jG
ol3bd5n+g6OUIlX+2JypCVOS9HnCHQWOQWyCK6Bwzxc+Ck/OxwZl6yNUSMRsnAZl
A2A4319I+iSVOxAfs7fw+MCKjm/xjA6TLzvdVo1Ya6rGbKf0/mwv1lVwMEsJlkN8
6tGLgf7mzCI0f0vVBd3Kg6FYcQYLDp6U6b7nP0z3TLhqIvMjj0f5LAkR3czAO9LU
oKFndcheX5QRDLaDp8owtqbvTK9oVVeQjdTcVKUhnWFHUQh9I7ufThN1UoZ1pw7s
aVKJ6fLucxcxqZ3waaLbS49fif7ZuscWIRspwWWSKRwR7lyYUH3NJU5iB7taGLle
8LamB1eUGfHT47+t+tB8qU63JUjeHaDJuhSFoQDmjbtloZHjMRomwGsNGKEI0gLI
I0zm6WG2dftVCn5ipLw7cWDD0VMmGfnVXRhKce12YRg1rm0WbjaaO+192in3olZj
jCf8dzcwpnwbQmr2CwwWUOCVB6aYLVub6lDNyUp3H53Fi6E6k6/RG84Aeh0qoGgq
rza1M332ePGJBBNdHdDC7Tgub09I/ELWmZvJicyJ74RA6tVhEdKnhLP+lfW4r0bp
JDG6FZzgYPCk3bnr+5IO2Z9/xzEp/K7yxtCb/RwiFxLDIXVDo71qgD/9RShLQs3Q
4hZvkSkxDftabJFuP38aKf0szmWyZ2TP+7VELg/DD2+iWpzaniX4nMCS/WhkOwIM
QF7PqG7O/3u+REWJH/sFp5OKLTBB6Jau9cGJ8L1k5+5ael0i8o5ZbOVIigHJFV1l
IED9INctmIlvByYjaKmi0bwxAX2my23fqa0Pqng22Q0WsrYoyaaJRxvaRmENsmIC
UKEFGFxH1MNoSFIIXflxSeE0I5EhNK7/QaFUH68Gf/zea7UL0AM5K1BfghvTDhvt
YKkOuZXrczAQ286qLiJzEfzDRk3LoPjrPLsG4MICkLNihvL30QnbVzXtwPJqRb1E
nTl/mgogsX1pW7TtUA/eLA56L324PaRZojLAdGDC78eoPQ+ZFelmT4UDSckrvo4O
uSglhLf+Gc/XangxMq4ZRARZvh8K9kzKN47DIOkvWRwPrDyCuBWlHiRfCbtosLlb
BFSH0wnnDGe9Wo2ISp09OjLuI7xQ1beJDS2+gYnn+PC8M0l6uGCj4fhkvXqAQ+pE
SqQIVJtOPORXhMFPFCud9i0GPHFMzRZ2dADIrvyZ3I4VO8vt9kcs7r7AqHlQDfum
dO9UHkRCXabNd2jNfA9E7t4PTihtsPdpf3Am5PtGwNsw8HYCYQuIPOnAzvpp2Rqe
yleKdsYSUQ/BP1QF37wl8jcYotILbDZv9tY3Utij5I0y9jpigN15ylCcfGx0XA5B
O5JpWy8BF6niBMPlYCrWMQRLVY5U3Zl2GuL93vaSiwaLlHySto2xT8CQQG2vEAeH
2G0IufQynwLTJ8l7Zb+NAr1PQU2cX9bgNbOUdjGYGH1pzGM5gBGyL1nFFn0hZwFY
yU4VNhz8bpv7Wx6LPNN3Yvwt58XCZeY3/Nl+tHsrYZqzOwHH9+l4lrf2WRr+tWmD
COINUHleJc2KbuSRDq6YPodzz5XXOY4XpQ9/+nQut/ahDEDMel5Vam8B48cPi6nN
WAXdAlnP5BRO0N6K4Cf1iwBiOiPovzJYwvthzR++sbzbS7ApT3X7nAqxVQNV8ufQ
h/hoSKjVLJliAAXimCGePDcj9Xik9BSzyU1yUDYY/CXq1r/8gbz+EZP9gSsr5fYk
KkWE67+p+3irnOOI7GwwAVpm+1INvMebA0DvpwfH1A5BLXzkXS7dFvT7Gt12mx2N
/gHVQAfnzCbRA+GR0IL8mptuMoznL47QZ1DJ5eFlNIFrjVe911fBkwVcLSilpsCf
7i6X8f2+ReaVFYAkdqoe9cT0B01z1onMu4RBO/8KvpEliqZ8+QJJdBCap1WnlOXM
dsTkXZVL3yVpZtHYdY4zOGLp1qomapvv+T6dEFpkAGWBXaGPeLlfbmrpsLBWdIhc
Sy/qxORJ3OJ4P8nnDe4HfyeMVTnWZdyCkIY/rnrTayK6Hka40T39AdtCwxpymWYO
ws0Fwo6RzhmC31SIfFiFfNIOS5/cUnpZBsgOs/62ks83AL+r2MIYXKdyA5TQuUaN
HrqVSTK+yCmdnH5yPQNuzoXqwL8HxerN8yOOeB2jZ6rgHWDpOpaL+9yhQUsoZ8k8
rlQ4BgB22QWWpTIDPuvU9NSzvulIv4W7+9Kh4ehJzMWJFUF+DqnVoVCdMwW2rPyN
XUqJxkzi1uIWMRY6sWeTb+4up2oVELO+RlinUmUsHlpY3JWtzKiH5A3LK6u9Bl4z
kr9rLXkwUktorwPwM3Hd6YBSJkgS/6UdPomCu+SM4c4vBawoOsNoAB9m0rePyhp6
NBXhZVAoBpW3sZTm3bqXXPFbDzYB/0UQ4dbJQRTNfl2J37+bG5f6BObP1vmyxQLZ
de9lZPw6bpHx+8F/daU3dqnnGHCDeCeDT8NjA44mnzFq0/gZJEwoGZo/wdQQzCUX
dt4OaAicstl2ui1ihn5CeGA2uKxAN4O5zhVSnqtNsyTlg80d5/KzbpH8r+YVawlO
Cl3+jrGjNzWXAUOftlOC4mr+byJ5Qa0TEo2quu1vigOvjCHz7gN5GmFKLjnN793z
xnxoneaR+mVdKExRUsDRlYRJrz165FlhfZUzeaOI/FOSo9qHNxvIwD0MAXcciZfa
3/c5mWIKkOEKVfPK3B0O4tlvZKMFA0unvL7NNgbqpKFb82Rg9SLk1qsg9ossLStC
+GYJSvyJW2Imug26ZVwdZUchwLqszBCLflvypB/dWsk2EcPHD9e0rS38pS2AgYV+
ZzkbKc66cLrkrnMA4f3mQvk3EyNwz1/bSGmsr+wrBS3zNPIe8Z15dEFrCsdH5tR1
CGwERLw44QgpVW72YsJwn5JglIiYKtwCpgjTkmKKG0pyzU0EX8Tb9alFkWOgGpI6
hhINDz4N40Pw8TOqZm0CMOi/hu6qQojsx3FkSiP2vt0jDCk1A6Y/9AW1EUJCPakE
iyAqhYYz7oQEY0z6Rc5UoHA9N9MEZerdI9hdqmMt5Y1EAu7iqeL+KJX60r8yUbGA
KTpAW4jaV86wVAP95QLYNkGJZxi6uhUjCRx6rXjlrIbDCEA4KV3shIyyrgGCJ6ml
aS+69HIESea7k+VZ+2zs3hTnSUD6rtPipQRrgrOpLkmB1dHAx9Vx2aZ1fCYt+mPi
xbm4uPRPXqhR9FoXXF9333QX2aar2EVg4oY/QsT4BYOXoKcA0GxRXmSs2Pq5EmwU
a0p4rvjm178kEoCc/iKnzPAhQOIKGoe+6nSbSPUerjHzL7gU+quOWtK7wbswwjTB
uHvNdm2gPWuXojcKPtjL7pEegsRO7gDwIzQBuvGn9F7ebc720fuz2BkMjWRVpONi
+T36pe6OnUAWhc+JNPtUhLBQQyoAARRXT2fXJ41TkS4UqDndDD8J9CmbmUuR5MmX
B56jYUM2WU+ozaVM5KSwocq6e3pDh6fSKphwEzH/mfKjf3LeBeXe8Tz5HPQUhjdn
DZzXCKHv38L9sjnUrL3zjL79V9wCQu/tufr643/KHEsrLXEXEchKHDt30QxXOEPy
5iC2dMlwUT6qJQXHX0hl7w==
`pragma protect end_protected
