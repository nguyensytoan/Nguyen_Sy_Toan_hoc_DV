// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
tQ8TAi66wCqoYiADV5vwC03EGe7W43miR1M0IWzoHHxOk7/I2WdevVUr06iPm44duwcNvhwrZJ6E
wPtoQDElhuPSfj0wKzG8R69OaoEyNYx1MABQ4XYf7v+vlELzPc3rLi0rD2nrNi5Z68WXbnk8yA9V
uv3JmK8RiTJ1uAU84ufnIW6xbRkIdVVDInVVUqm1az6xF2TKUax+zfDx8tFHsdT1ILS5nT9pA563
UiKFf/Pr1K9GqC4GMHypcigq6EgwCssMPTyQLESLu9ISsjk9+zG7N1ByBFfNx6Q9voaqfZKlRbdD
tHMequE+Z3DDwzhXoptFBmieiSC/tRwSKaf45Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 12160)
sBq14P9lEABiONzHlS7QVIKMiA9QTtAUA+ORIiWghgp5qkGW2MbPtEAw0LkahD7LwTe7Gkgs5K+X
mJURCtGinAvo2BlC6VBvTlRA6ICkJx8sqtsTvPCBnplX34SOdP01ZW8m0XZBwCnkorSfi+9LKpMU
0DvP1JR7oAsF45gg1xCRa3KUOsbUUE3cTyAo5qEhMMJtcByslQLJosO+POp6frRe4Xzy/ba5pyhq
k9Fclp3LWxUbc50SJOuW5lDp8mKrxrqrhi63+eMsAW2BK0PgMeJYQG0CrPaXBr5HYDV7g6HHFNG3
7Qrhc/t4Pr1dGSFI76bpKOuPWbHsqvr9StA8EGw8yOZFnJrNor8G92SxVM3fpVo3MxT75wLamMld
YX3/nFJbYH3E+WuRdOJYdrfdZpYDSsEtbiwwSXx51+aKY1foA25ecGtsjKYb4l/cFTm45NHBWzee
hN0SF5P/ya371uU2VD62oEujHmMuzMGcOgVKhPuHRB1Ztn9z1ySCDHnD3BL4KFqYgHry1PX6UDVz
IdcH1F8nPwRHAGbPI5eLvOxc+wyNG8ZK/6J6RGDavPKMJPXwXpwEWcJFI1/SCA7kwcv/u4BCMVB0
hFELUUrF/zdHjhDywqEVkQXGcv8KH5fR5MUXhrd1Qx179bPK8w1MHxn7GsawMW76fA1zQnLq8u/T
mgMJTe7WRc+8CAa4faUprjryEpMmXfgNePchkx1xmFEDZtKIXO127E1YPwgJDoEn2eRZuI+3T7Wx
e9pem3Ieal/tEXYyjo6+RRcyXj1xghiM0F+ORezYMZHuykLTBYwhOV2F0UUKEtht2EQ7PjhOP3hb
hr5mw3Qtms0WReeJI4iDVbFpR5/DckcSYae8njbLvQ9FZuyDY37QJInEC+0c0SsJD790Kl3mMXf4
MbwU885U2/MngiJ5LRZiP1S3fM1HHMNGIB4eM9RJYs1Wr+b7k6Xw8EZCmxylpXwCQaNgpEOkNRNA
C3Sy/HOndhipPmWaB/wlD64RjtRlW0YCsOfF7lvjfneiV6yl49+9q61zUhVt4kVL2NgC4D6NjcW5
BItXjypOdSNyVL54yE9Zs9qVoK/A+TbscNRwVZJb90ZA2tl4eRpDS4F2RJ4YzAyCgeNd19QzwYBo
UF3n3Yo8asHeMrzu8Nlt8glglJTu1oCeCq3IASnBPWbaCHu23qkA8he6BMjgZeX3j46bLsy9DoUh
Yg5prmp8yPwm37hIsouMvx2PvykYbztRvW66KHsq0Ph95j7aEAM3Y2wSEE5D4Om5QlkUB9fLZTQ1
CLhyxKt7fgBHeWXqSqRIzu7rnU+PsmcYNlFMPJcvvsg8mZPCDshGnJHlAiOOWglMhyjICWWIb8uS
4YXEYP0ueH/bMekURl1QVJq/IEEO30O9ZQZae4bQ7j9EXirqmQHJzriO4WlVRYtt9BpHGdtFnNEc
R5VX6XjrX15loaXZOk3h7GkekmRZO9YY94wMFZn3jpNtolvSAvEpDfDm44mdUiApHY8GcLLCWRUC
HBhwffH2kLY7JEwGWKBRBPKTcVJ4nrzS/SrdJrcnpKElj2AsxrlekbaAab1XzMl6NQyyGush520E
lyie7E90F4uRpsjw1qe18EaQTKHiE7ZDiaJjiO4WDeTAkR0aaM/6YRGg0cg3l4nHUy/x3uIUgnXR
EX132qPG3zGvUaHLdWkbKXqSMP7T5CXqOlLtBYCPSqHaw2PbiyrffVPCWojlw2KboVMVqO/8NUKZ
h43tX+vQ9OScKjkd5yE+ETl9p/u+Hwi4A9kmok5v1R6GOz9Pd2eP5aKsypUnOgoZtpkLjwZX64pj
5593bpBjueKxzyUvCfjw5k71n8678nI9ieSoQwD0x+P8wP8Qtwye93eAlk7rIQg1x6Mhz99fJtJD
xnAICMW2z4+2qS/k+U9X9SgZn6F6c88Nk/8cqbATCbDC6DjEEXZFbbyLQqa1kRKWqhH/vT/HSYcB
YzP28zd5BmNcE8uf+snaCKpeavQvXlSfBr8ovW9WCJ7pd+rfxKVoY26OzKkAnWHn9Eu0J1e8yvoP
BHAAdUFe9rEXrU/szrXxDu2ofDUp8OMewigSjd+CS1NlfID2X/3jCQJNIWT2dPmkNHObUPfbWXUm
y60314VlYoAw4wmdHpHy2ZrhiNwtb6pLtHfQWccjtpHSlbpK+p4XY6VqjGKNzsTdXrR2zvoAWuOS
gj8wOFyKvtlpwVVgEPcJal8jUZelTB7mOZbnRRMcDlnP8VMxE+qJ8GXojEOnpQcvj34Qdz8XwHh+
7gPItC3QLlqE9KRW3mOjB1CtJ9iTvzrHaSyToj96GF6fzGDWPrsNFQL/HGLuyzyUVoZFN5GmzMSP
UqOCgaANrGdxfaBB9Jk9n1oUcz8TygPtFebk+yNuuGYKX7q5MKi3j3XPLva4A4HdSp7OxKhbSFcK
cpI4pn49JStciuMjDfbUcZur/qIrbbJEnzsaXCmAIQQpR1HlS+77KoWRsHm5oSHbmZW8yoARmQ0O
agO0xFdRjpXGFoI25BfZDKJBXpeDqBGfeLLUjr4xstHXPqQqun4nP4Z72R/AUXMK7gJEa9U9joC+
hD8x9tGWvTYYFJKswuTDyJTJih8hZkNkT0MCGZAYsUynQerVu3ffJ61K+MOiltRdsEbQnqhZ8kqN
7vKH2hyT4ze3Dy43a7vejEkvzbR1FAJeEKHbFc6DT/Kmkg94AR53s7PhZtbw/kzq73GAFU6pGHbF
lPSuv56O7txX5KXIWQtQu2ygER9q0KTXrbeB3M/Z3ywZGvPaOTuL/oGPBgSPNel87r/FXiVBPeOP
OKmBzFWax/rjETHLc67+Xbd3J99RQQouJuxmmOzVoBanqy2qLmU5gHRsXKDauf6qvglwYdbVer+y
FGOcAfaFu/2LgDq1GFlXDNyqkXjkiCKJM65Kr/bDsh8a7CXwolv1QSLWGM1/fJX0QOK9dd7XF7Uk
vIkoJMMe0ie5Hj8XAimH3al6OF5MBK6pRX7QjxC3mDw+o1dotTi5e8KcU1KY7zLWgjolQnUGpPS+
eIZ0e8C5r/u/SEgVq3e0VELSHJw9BrDkPYh+xwyDKOt2nvzDyI0NCcUfI3BAk8mlCgbFeAqLMpcf
7MBOB+t76U4XxW46+D0UAGoWlWMxvK/Th0kMHzWDo7sVxOwijnDg23D1M5++JISRigKa/YL/wvur
NBh8kyUvGsA9ym6ysMLG6s7bsBItFTx1xIVIRtKTa+l+nfNkDvrCnEEPtC0CUXr4CH8PoEMb49xu
RsVJeKALwCCLLgM/glmSeNfNDDVl229TdkbvDIbtcll5lc/tWVSiUIygHuaNpZSPCa/lQ1Pwxyt+
xrUzilaDMFBzeKaJkxeLqYvqFJysvra8Fm+d3IBlXsQ1fxlap+EXTGNyQURRrIAv74JrDC6LZgUg
yByrPkwk/IxI8q8MH1PvgCruUhb/S13xrYxce/LjjyHIXkgr/8updUyz4qxD6hrwrIDPXbgXTBcH
FO+rqH0tee8xIQ1NIg3ogrNAXCUxHZctKwiq/fS3ungwlhpYKGjFpvcPZA6c9XvbmyVVqWfZE1an
kztG91PH2BjYkQYcPm+BWOck8x/HQkORPHHKNtIla+56ux0JZ5zeJs2oBfO4z2JgUUxBQ0tfpEsN
4C8Hn4YK4IdniB8PV1kZp05Nnai+wtu26tOu7uPwcBd0iV19CJYGDll3+hiY7n2a217xurZHWJw+
dttioz0onMim9sAwaph57KIFC2X4AgXY3epjbpX24cbdoqtLQuH5iF969UnmfV0XaSdtbr0Tnii/
jncoMKnnW/JU6D3+b5NUchXAONUoPLXitn85mrB2KxvcOYYssC6uACYlnKTxQALaprP6SwFyXI6Y
VB5uuxfE6WBl4pIuQVFBpwk7jL7559s3pQXWZppbbzTVIJj7SVxXqZgD1yowOku4+iqxIyETD08V
kBZ3Y1O0V4NHz0nHbhq6hq2vR1EN8OJi34xx3FzAZEgCJ42tvZUJ+VhfXieEkWQy6zadgeE7hIO4
trsqDz0Ng6Rrvn/hShtmXGYhh6TVJptkNXrf+rxYPm35N5+45vHoSeo5w/W0oqIRRVQDPXXS2mL7
1Jqlqra6UFJ9WmppbSQu9GKI2ff7h7PmXdOfzrl4iBvHtAtTj7f/zFH2bikAuMB1kxLK4g60B9xK
e9Qz61hK+lDHEPnFWIv+sfQBol9Lh5LJ5TVr1aylCq2tcFXhtQ2Sxs3ZqMbRw6ZTraUHgKIO2X8G
nK0GrFxhQH3Sz2JM7yt/6XMlskVW//Ra10q3jUa5mpeRz8fAsiSmlPxDyBwJkn5FXk+cSuX2L+Tf
KyYuJDdD2EKwwxYwcwlGRSxgS9V09qVB1f83GeZ8/KIHRp9obN7wmYPpbEaVxZfqClYAf5AIufPt
gGu7IcEVTgs/wxOMvz08Z4e3oLrAJqkWPqZ9/XF2VqcVOm5Av84M49htjtyesZMcml7EVzl9dB4X
/VEVcGI9Pj4btQvUus+cNbBAre40oP6MRB3x5w/5ZNBuxAaLI989z0n7t8QA0AeSPPXmbwNh0c+p
lrVQC80BuQqv1to2dV6Osq3DQLUqdc985W0cqNbpzDmrbSKrTgAjJPnDOPrGc0dKqYLYwt+NnRAy
Zvh/Hy9OZVORjaP56UhRLOF5zpSqVRaksoQYe1cbTsZi4ZrnNavE6yDvn1jXJCmVuWemdzXC4Icf
jPx8XKoI3/fPMfUB9NhRakFFpqkzzwagjWcno78B5JE5C5kaZ29NucfoyRYQVmLHPVVysJYmGUFs
0T/gNPYaqqJ7IvhMHq/T3PBPH+SpdD8IUIoQH8ITgrp1jdBlfadrweNGVkTuj83MJjaqEASR4FkW
KVcEfO+8nWhl6ekVGlheQb7uNMOFgnoI+5z5PY1wFyVMInq5SH/DhnG6+GgRZcnJZtrMREnDnoDd
KNuW9kSuuejMFd40mTCTnn/GUbJ+cMdPF9D3Kiy7iIiZx7uHDIEMT9J1iyYhHhGumAooZy/4ryL9
Ris0l4jxVPgiq3dmc20c3OBVhba9Y4jOfoSy5ie6yHUT+1q2JXxmAZ6/ejrd5lXEAP0rKi/Vnr/R
v92Cpq58grJKKkSA51R3rjlVhOB+MPfPEb6c3T4l/CfaLTrYSQ37/3DOYiGkG5KeVJ+Dfvc0EW9A
7Z8i55YUEcTZN+VGGxdtpjfjR/Ef6EULp8cY4+rgvUCkf0x9eQi3CArnhO7DXnigdRM8lIn4aDf7
C3j3t4aqW7FUa74UwHUDoFxKlvp9Ijdd4SP2zdlQDgLWpq0I94jIAEoFbZk8Kc2rg6IHD01adZfK
i6k+HtrIXhGVlmLJjZCyRWnzw4iDFQwEOLMtK/RXvAN5Kk9HCRvlPze3oW0ypDHu4+klOSS8V3Ea
+bcmOKQqGkfwJY30b7ywN9aHJGh5G8Vtq6W7I9ys9KnhCrbzMITZC/KnFr/VD5NE+RR4KEL2pg6M
56Z5E9Z6H14Mxq+7507rIeKqeTQnOUflyKHl82n2f7LgaPp9HJOZ1Hr/+5UOKmh0YN/qyxuekGUx
9AhD+6lydwXOHkiWwFUeT1SEH46zNehyBvYtDXSV76MX4NZTTT/m9+MmZQ8ZxLK6pwxJOAWUnBME
/907WRkX/s6TFpVEUgjKYVgV3dr+z7cbmNoKexHE5By65X4EdwYXZ7Xy15cS/jjaPkfpy0ub001S
EcEkXT+0tehqf3j4KY0/Ey4TgEnrCBwG3HcHPUrRY3PvTOqem3JE5rrU2YgVZTRXgA9vVk1qUyR0
y7NjPiVXkRHpTd8glB6ZpiZ5tUU2qvbC1Y9ub7wUao2rm2oEeK6ZsYquZjSyoZsXcbIT4gOccvFh
zrEpSyyAbsZU8nvxles3x6qHubUablWCX0OUslW8UjWNU1fAXhPQMu+l/u3ulMwufj8zWPtI70J3
Cu2vtwo4/zelh+tJ0yZl94JYdp5/37QiRNl0QpIu+0aGbHmr4+5dhmTJJT0ZCShKd9HHpM2oXT5Z
wzEHS8Jkw6ofQ2NI3TsgOnchRbgFnAp6TVhvUGAmf7BAVYV974PPStd4Fikk0tuFIw5a3qViUWar
jxC6U7rl3OfHeesgW8u+7MNbteVX2vm+OfgRBDDA1cBqzFqmSGKq/61g12QR37DMEit7E6fLfPFt
Lh/g8te5K4irtVSuqvZoHtLaUhVGnrSwPTQ785gwfyreUFyopff3A9vv7swtVdH/AwXHshfq2EbI
XSp+wPnssT5fo5CmST3cKlxXb4C6Pwvxjr+mD1xDoX4iZgvYbToM3h6/ZS0aGqoET7/tOrC0UuM2
OCsyw+3bLXSkvtg1G+EwUgKntORldvVrxXEQtg75vCA1lcs28TLOl3OFVLPIcS1INICPqB96/6as
E7uVKFJBeG64ZcsB3RZPksiyMzMXKi1tsDInFiVCAls0WBy5xXIPfiVWQT1nh4q+ovTi2oy//KU5
SnCImwzWG1IIP/xBuPQHM0Zcsqy97gmTO+KHvrL0uzjBaD893O7jH+y8Z6Y7+mTY1rnlglRgp7KT
ilvY2EWtA1cbxD5cr6o6+gIS8Hu+ChetIXIN0m+Tds7hRlxrB6/0RuEc2wt6OD5g0R6Ur9NmNYGk
QPH99GTUPi9B4qs0QKdzDlDNJP2CrGj1D5NdSswBEeJr9H6zCxBB9MCzKklMp5vKfnJVNopbQZ0j
JMmQ0CBGjEYdVibBEQnFCBKO4RCLIuBQhPIKeUR0GlBFLsn9aPoHDedbaXYBi/jMtTgvEr6Yugbm
U2lx1OG8DJlpdhOA5IyhlxNxNKKPmPjD7E2/BzztLDmqQqmdyG566Kj6yktrGg6STa0AnW9MbDhc
4Iyi3nd0ZQmZGFGhPi0HpG/XOul7Fm450e9W5OoflH03VDdTbItZ5S5bIk72sShuYU6uLjqArvOO
BQ4cULCZR/8ani7Dx8XfvPEl+gFUpXQn0JuBY7Kkw+PvL11uA5z4mwJ7RJjYtYs/GSfCqbO7Mztc
zn3AFINQbjeF9xR7MaQ18vI9rqo6//bx9hIGZS96n8f45rdb4+NyT/ZzB2XqpDDwls9KDDG4DY8h
DvP2S8KEHAAOM3ApV9HlwR8cjUx5VoLv7QVmbJ44yQ5f4GHipxkqp/C+LmrokKMgHL8yX98z+Vab
lr1eNv1/lVfm+XVgtddL9GF+jV6z0XnSVglZ7fWvyCqomga4VUTdvC9t03eAWyuy2coQPWWSRTck
gWvDUmGI4GRLgUVAIVwhyMqB1vmTFjQIzQ/TUZz5IcPDqDsds7JnLBEIjUPCA6dTjFrhcwB6vlYV
2UdEbdzN+u+ngC2d6sFdEqxE9sE9YjKCASI3dWFU+VrLmA6Y6ukVYF/vdPE7gmu4O5cAME3EbjuI
uiPk80LWG8JPeRKGHTXccpuPM/UUoU2aEUWA/P+raHmFbe8jqDw2YGxQG6IVJgFwf0q53qzqB60L
pK0LZpQiL0WwFdbdEs7jYvTbHP4XZd6GKV4mD92eUQpwoUYjZ05pYl+xzKHy2/VGDkZ2YmWFXbrS
8PsxYKS92NskqvjFeYRpU+EuVcyqwD9mlDNghpILPQOaZRhhCmFc4E/5qOOIBmdHKMlK1BIYbUZb
pW6yQi5EiHLuVyVIeiOqTm+CAdk9ClOa7FUnb/gWCZeIBW9HXrJBRFbi/mjgmtI/Ezg+bjmcZORw
bNklkrxZXa3KnzNcAVxRV5JbjgURQjYV+rGxV3johamFc5y6wUTgmcdfTUBefp7hQbR2o3+SUZ2S
AOmlsf8MsIwVIX3fkcVJE3CD6l+ITooMMTdkAz8Qefu/q7Ndl+I1TuXfWSWdcbOHXA5F7bbv/srf
F8Xi1eZaGBYf5uNXuGkwGYM6CEqa0WuUiMBmhLmLM2qxgHiXk2CYdRfogixiS7zVd4BRCSGsXwdJ
q2k5oNOrXKVdE1lGmtp6GmHwZu4cfZ2JxJg4Rb+j6F4P740lxhKmhheUkc0VK0z9LSCCQtbmYsur
ODAD1YQIGpR+GkOwKi0PuRsinEopX3U22lTqkMIgrgGI+yZb8lGUP5s7I600On5dL+vzXcYo7CD7
m5ypwNBPy+uGQ51hlmqpGCE8T8y5fZglfHdBxdndGkbKoDaUM50nLgQETsIZlgm9EeBDtEVadJ2i
+mlaR29wYlrQALBV7CfW5RdpTzyv5flKURQCyLdqUVDDoMgnpi4kQbFkezj5Okx7qPmnOxVbP2Sn
ULZUCOA3ENNDN4+w5jdm0XL/4ggADjMx4OwSOyn/RuQ+EfH9wfzT54PWwjDyK7Hk1vuvDiJ9AR5O
yjTfA7ttTeohxtD+pP7yJousrBXHqzl1bMKkdc9dAfXI+PzOkY3LizJpnXFF6vUPaoPEaTfFPulC
iTirijxn11NzijP60qUYuEPfPGrSHrW9dCeMRE19c0ZOyGjtxtV2wiEgVFYvwmMbrArFB3MLJ44+
jqGCB10k29ODgPj1DUujmDfyoaUmH9Xsd6gc/Uf10y9L9lfvu8Md0xt1EPQalQ6B+WQ/c9x4DEIw
lgHcsz1o/rzVTF90NK8zJnC3f+EjN6FhHHEA0tsCZA7wG1XVg+ql/X2esxBfRlvox4zu6ZH552Ax
VmyriNzLmNfzxkdjjjseM7q9kcjXScsEa34rKU6QjOJ8j3mzRd0EkwoIs3kV2wHbDtmYDo/5gMIz
p2LPvDT2LSxb2k9vKAXIiwoGkS76oh802oDZ/sbJTnalzRBmSwP8WxBfRNIT1VrGlznu01G/Z366
+nx8JgMsP4dH6rwngOVelMsYRqnacwCEQ0yvZZE+x0QkI6SDNiQR92Ik6x+GdDzMWW/iRPhH/QzB
9H9L+EdXh6DLW+i/a1T0HMpjsjJ3Gr7grZE/Td+4GM4rdi5GEnDz6XmK9vmR8FsoL3pB+HkO9OMk
vWDjP5/nO2d6BDX0vj/LNx5QHPjxS0Q8KsxkuTXK5/scfVeCc7/U2mrcPQ7jDyeMzRtmoynGo2yh
ZwF5Z0esNWvYmnFjA0jwS+YndEfK2neHBq3ec3I0K28VbTW2FrqJ7XljloSbjCdZ9F4aSVIMAw00
20Kcfvb+dHXgWa1lZ5onNFClA+ek/QUYctuSF3+hLLBnMZKZjXXVWSK2CLOfaOGmur1YhTQLtiUz
2T0Eyyavza6VE6SGuXKyfa+5NaQ8MKxMPoZImcxtcUhQgkb9dd8rdirDULWfVhrmJb19mq98LblT
GOdkatjj6vmus32wBKo5XrkrRvgkDOk5dQY9beEzlyEsDeXkvp8A8k5p7ZKLsEsK7YJrFI15U9H3
NgotWg9U/PXGOUTDEA8G0wVdDYogPnmr1Y1mHrXz4pVy1sLRPJMZmDOmolXdJEslxQJoy1lTmkzc
SO5VIf27cxpwe3+Yx1CWT472IljqVJMRiby2pRvbt/Fm9gUCZ0zmSdTxoYKPjZV5CBGd4EcAtT9H
1EK4qmCncpaXQU64fAI9Y6mM4mbQ2403yIiK5XA2bvoshbEBCyAT3C6hemIXw200eM/jPDAuUZxY
vMqyhTlmQRfIlCxIhUqK+Ki2IasSIXRq0IHBqJRxjPDXJYk6DMLHZDzBc9MM3Fka26FryFcSWTMH
PA4btsyyGZN4+XiA8Frmotc44kYUo1L1SEvZhNPaILBK1BRw49DS9b/t33l45tpnrxZYfv0bnPjw
cwn5afTh38hnxRaZ8hQSVEYm2JqMaf8LKToOo/kK+MeDLUKAyq5w8UoGgmbPA+zB+8kKj8YfG6au
rjqsPepMsd24gzBS4iM1z+5m0C9Dk9EHFVuGtHH8KEoM0j0B8Cf2fi/sc2EZnT7lvo86f3FF9+1D
jl3J/yGLCbFsr75If2RClDVDDp7A6ycLDfI2uAVuSaXsg06FjIhq9mnRy8ADFgnPjLowMjgqDy/r
oaF6/5fKM6b6ApBA25TE1aA/R9MBvoXJsWkARhz7tYiFJ++wPAOp0Qmgfwm+6hXpwSatXtPEd9k/
njsFQuhYYPZTwkFpW3TRZMTu7evdwSI7e0dNylBi4zEnvgrsTk+Txfx8cZwqUE6SLNdgsHp3VlEe
NWwyAuvgmXmStxgaQEyvYXTJf3QYtjBiMwo709x5qWrhd+Z1nwKveHRImzW5MlkKOYxENE39oZ3p
Nu7f4U0mP5E3bjrAHp5chM+NV2+q+xzXjGw2tycMLnqcYF3s/k4do1RoyBj7/09w4vs1BK7QF2gA
D1OJyhN8BgKd7YQSKNQXO4wJ53kJVKWXkH64A7K0w7SiUQEfACc26K/s8vZBm6/+KJwoHKzXZdQB
NwJq3kraRlbHDzY+5OC7rGqAc9juZK4u0h1Rb1x+A7Y3Zzdm7iAlj3th56wtzYmUg6Qsd1VBgT12
01vzKKmbj0oFHjh/HETEhTz0bBmJkdHph/nl/Pc4EWZ4zwOoqurZHo1yErUiwIV+UWvo8bzddRuJ
B3kjtuUkD5V/3z/ABfLcWMtBgZRQX8wOwxAZ6vnz2uyh1NJavHuOGJnE9kj8V+QhexKmAtRUqXxZ
ftRucQqiTezCR4pIu3VNsbxP5LkM3dSNpcBwPb1GLNUkSQKiEhMyAnhm5aOfexO7me0FnI5ltQoz
obfsWpidlL35lCnVl+Y8X8uMPIUFHjpyFrcSTpGWcV9DUirzeZaxpSSuqfX3VLBJ7+P2miEg02WN
l6Dw7hbFIh5WdJxI3zWgEUfNQjuGkZDyML9ZTs0UD4iXg4Nn5LfNCnUQrwPHnnZVwSlxS8NiolvM
nJX5qUVUFSuGxHpnDba/yjHPM8XJhOmSn9nYa2Xe4+/4et5KC0wJCjRQ3vk4+5l7gY1nBL2slY3y
JFwp5K4kgYTcCkI6l9FUMu6hcVAYofOjm18Hc/OhgclHD2V1dAhuefSxURzTyGCm85P/BxCEqtBZ
tq1aA5IMH1jRhFziGAcSoNK0JDze2N03sRMbQZTocRdKYBF41uVIoshMXFXBzeCCd0k8yTzfxCGA
6SCo96OcJXW2Wr18q3mJbexAMgoWSmObjoPs4j2pam25gqgwJLSZy6X/hJiUgnWnVbEio7vGJd09
7aUqQA29cN73PX3L3Wlf2cUS6Z/hQFLxvXupB08aWeJ8PAdwksq8K2ZecdvYbtgWLCEaV8yMesbB
goRQKVvs/vY4oaGPn1HJf9kmM26x3paW/BgerSLrGRzim5XOOGvNiiRrhPhI1Ea6dVEU3BNE6xRW
4vF8ee/5Q3r6Tl59eqGgpItHk5pbiiBZsNyZcIIr+anT3KPjl1RSpZHlIYR4uF/agy5si66f4gaT
OA5QSaEb3uQW8Fr4JjREYeMdzLavIsDhSGhn2j3doKomD53UtKJ8v446d9yfM+4f5fzedXuByzi3
eFkvTTRZIvEJwjc7Nu79fkN+MVkvQHMQ7qb0RLKUt7JTXNW877QdcA4LcOUpWXTW4rT1yMOXIHED
Mk5Nf8GQ5n792cXkPyCQ+jSts4GdQ/KkiJN924QOwel5C0kvr9uJSgrOzXEn5299JHBtGgtvCKYL
ZnZr4Hyg/m8ZgPWeMv7YVpIM5PmgKdx3efdmD5sngbGqPpwNEhPXY687cZCnVe1EWv4+nX9JZ/zI
LfIwSowDB9kpc2Um201T3H3Y3fpRa0kH3Lu0dv5YCrQLKUhCacl+X0UZ36q5gVOibH7/Rjm1AE4y
y9RvNPVSkWRUkgEQ3yXVJ+7vyr12MwHvk9rtnIF+xQo4FhiS0IIzpmCDsUxFkkGv2ufRVzkjJUD8
fL7cfUf2atmziyVAygbbi2uiCY247QK2hXBM6U2aZs4FkRlYwcnt2AeIb3IWxe3uJJjmN66r7cTN
Icivtfiu1h7Ok1k62I/w1yyXR/Q3xLr+PVUwILTYE4bkSUjt7oPzJFjRjbdq14eTaGvt8QCIDyKz
dApNk8ZWY/gGnLAm54aqjaOFDInu9dOezZTpjsmt7p10lVgeY4ctHAb+i7RCtx7HocHn3k+qCoku
0GmkIIse3DrgEWG6BuA8ogD8QE8E8mVBvGvD1I3cr27rfHHEHikWPRLom45cdkctxlvG7u7UtPc1
8KqvWOlQsma0/YzhvDyTmEr14Hh4kqUSAW8rS+22N0x85LiLFivfKbdoBhdQkGDHl18w1H2diiRs
pkR6uaAeBaI558SsDeTt495/xrO2nD3fUxD2iHaWPtoB1MPUBFe6/57yWggJfF5Aq/i4gkKMaef2
CDhmvfhhmmwx8dioAfHjPiR4+prdhb8NV3n9sX/Uvi8HJY+UEjVovaJunKYPYxrdiPNkmjfkCkoe
jRImD1e2WfFALWmQjrkMzubmKioXWW7LM/blYi6wFnkbXS/TyC8LN3mJYn+HkryP5xy+JW43opdq
r97PFkMPcnvR0dYedFUgmM2BL/pLONyJyuaA4LZL6a+U1QQJa0mYQtqRm6mDWx1P0MH2Xr80WnhK
C+wf9fhfaEPeGildYlzvqWRnJndWA7fbapNwOzY6u67SAe0iVQtmznInmq6FXwVZZSE40XA2SKfo
3L7EXlWXCil9zfY4bBaSNxUiUzW7ZXAv9YEUGAJ00LCfOmRoR0f/IxMWNX5fwAoT0Ymoc+YDW/zz
DGJuZJkyas3uQGrQcRtvE574B3eCx1NPqsAoTka9R/x/zyNGKQ03zVBvTrf0LWvBNAiwlqxxys1F
qzqLO29CX9KTV3kWVyjPu1xjUJttMXjmoff7yz/BL/Osgik/OVoV3TQquUF9NDyZbm4uI64kLhby
op/W3Ll7vRVPDDily9h8D3uNW98VrEZg8/oy+0F/AbSJmnieH8PBJRrsM1078t4pvXeGh4cN8aRB
IJqd9YLNxrKlHO/wYdEpTyyir/3amP+PBn53KZBZY5eY0ET65z0ELinWB2dIpvZf1Xq5PIV9DgGJ
BHItjrBSVVnnZI5hZ6JpYK9tfP8dg9w2uC07xVnG+gxAuMMZme0IwKa9bJ2Jp3Cy6ULZHHFN8kAs
TWcGEBCoeV/f+nsPY9S/WXohaKk8Ek9dGBa60uxnXOaaz1Wdt4n7XFjRsasYqz8aC5eNYBtRfvLG
PLCpY8GHW55VKx0g/ZlTomldd3yhI+ke4eniue8hIYAgEtoNWZ6xtxPgRneCcUCxT6iANMdvvxE4
aBzqLNtK92v3W5rtIVXGCpoghDCioYlXMjeZqNwYUKkCU8Jk9rlRkYF+JGQZ/x+6t38IExS+bk38
g0NSWjgpSw+ODlaxwXyi+J1tDFu992YE6IuHwoxGZE2dtmqDW9l2XGhC6io/i2pwEAB+Hisx082H
xABz8DnGMiNv4zI8628UUiSeSEBuMxoycw7o9d0W0PZbQXG+jtM2kusUwRcx1ZCYspkdZtnh8daW
QR6naAnHsKnw6/oYS/LJVGtFKXNJtMWPLBGIG9MS92zSkspeaIQ8uS3bxlAWNo3YubZbzgz5WIR2
i+WaMbk3yXK35vHpeKqXa83tU1WUEYG92TvzQw7isLs7dfifZslv+usrmhvJ/hiNhmj+2tmrQN9U
f1gtRPHOxWUSxlOHoCLGJVv7s5DqrqJ+eV5wStA8mEEpK9bPe51+lRw+K4dk2T2mNgm7Y3xesIFH
ZgCAwm7Mlv5A4zrK3kOQ+5gvERuxzxby8RSuRW+HxQbld0eMdeSwUEkMlZ+tmWiBOnG5XM8pSlI/
FAESFmsbCKZyCdO5ZfuDjERjulAtNAZkBOCDG3lnUnwsU7k65lSyQC+8N9SZmy4SZE6suem1nQDT
XasU7F14F4c8W4kuIJ1zcYRHk2gSF/FDx4qBsvMyjc9348jxVNFFnxwnDXLpGmhcV/FiFk2fJCL9
2cso+Dw+/QTjsNsADOtDD/vdFtgxFcIU4W+JILWnNOWc4QyhpiTFPiKl/LLQ8EXzwGMUtyjTE35d
1FKsIEwEda2vvR7MLsQPGUbJ2fjSQB/AiuoZ0LRMt+r0+4172g2ImwdV1zuvbsQuvSCNn+zzF0Uz
/Dy8yqYtY7x6hXkOuay8QZqtr9xTr9ZNDA3kmj7Qzbn+RKwyWdboENAFpafYLkXzjOCD5iPbhokr
vKrW+ccGErDd59mDqhzuI7AZ0e+ikl7ALtoeK6F8fq5nmY7ibl/wth1P6FZR7lEHrtog8T03INDn
eS0EIT1tzkkdTnbr8J3XakBWTHb5yNrUbhXs1evj1fx/vEQ3TPiXHRdr1YmowGl92vC9aqg72cZo
mH9QVU2MN2C4OErXgySFCnn2G//DesmhV3q6kyhFgFCrD4sCSvJXe44h4m4CSyCHJeb3m3gZlVVo
1JrLVnIPsCzMVmC0Oq9H7NVRQ9hZEaA8JiXt6S4tdKwAQZfYtPsIdRQpTzgd6PMhNQQMs8TqaxwB
vs3MlQr5t5cezBGKKzuojSBV87fVILm84KFGQUSdHoVNNgiXuPaKFs4CCRv2Qjnt7MK2iyUNBUFV
SdtD0gsPMXjaw8RSPcJtQBMVzub7k7rGeDddIJ07tndHRTwTwglfI91ZsILuxUyGUqboBgcEjtAk
1jY4odzd9Z+IzOCnREhxrdKXC7iTEPMHo1k5ngMHoybfg5BJEK+1pchXiX8/LCt8Ntwne318Su2i
z3b19g/1ojWf/ducYmcFWjWV2rZujipgNDtmbAM1j496ANTzMhW3VXffz3QbGvT6+872c82xZp67
bZzrVu/aBFANfAxjqwe94/XwQQ4+E+0Ad2nW/Vtvw5/HFGAx276mDRba0M1n8zO9k9eJdsPhb8FR
1c9L+Vqv7nis+PSBrXAQMbwdVkinOtnDM1c3VKgVcUMVVwgQT/F0mzdijR3bo0PtEZIfz3nRB2+B
Qo0STsvTRNtGTTTF36fG5XgnbZ97ACkZOc9ARus3roWf7yYEFIpewCgO8gAOdRherat4LPQwF+iA
b2sG9FtpUHiK5a+YMDV0EPVN9doxDFhDaszGHN6Cnw1epbmf0aWwcof1NzXkfQ//PGYribFvv9V4
GjN3SdUdXvinNPUhjn25kt0aMEk4wyS98gSOVNXEZcSO5QbM+M0F2/88qyVxTnOmCku8snGDsRGO
KmabUGK27zOPPVbCqsstaacVKcPWcmhdMNwqf+Xnx0uzgFNAeoXw8NVUVPcgV5jvy6DoMq5uI6qZ
NLbdZkg/QLG3QMZK7FQeTG+a/YYd2PMdSlSFdSmGPnWefXLhD06lmQ401qKoCrmKAP09hCQzCR50
0bnsARauZy5iBkhJVvxaxAA0wxADAYQufGajRGXXKrLCv/etIMEzenMTADwSq6h9RPscF1f2/XiU
YGJJSq1X6n8xR7cARY81QWZDdKTekftEJVyncwtV3ekQrXjffRlDJgMs87hZxo4pwBqWB7fWcQ4D
cylTrMNrrCdjX5Lm3ZdEi2EMimFQ9xaxvpMmvIIDOfX3ih9KvQzAcW1VqtV+y6HiGYAJlu9+eAcd
eEVvjydbk78Y1hfr9GfBxQQxky2tJ7kYcfaiJ6PhtJPdiHWD4CsiCl97Gn5JEOobGPk5MKy+LwK+
QimRmszEnCw0oR6JSF7V/ABpImcwKAMl2IZs1v6QQKPcvI93cwEZrNqnlkmFD+DHxDp2rKHq9eya
YLUhdyw6bdBUWD3HP0+c1559bDpNt8TQDt/bcccrA7XgXyIFTy9rMIOo0zEHLw4GAcX0/I+SVrtu
xCMkDwDflvfpjreGk42AGjfqQ/+0KbfeMXvPoM2Kd/xdWAeHl34a43JT3Xn+ThfMRgxCWM71b8m/
HC8hs+1jiwQ13SLizAml+rylxzEFVcPezIjIuqJXLtMl0mfwipXcORIHBaTOX7SWqPdFCjIhGQnD
4i2xfBLz5dEVUzv0IZb84MWQFDsxfXq4wIkiImegHhtheLomnrxWskHuS0fZJab3c8ZMtGTA4svd
ArV6RXZeU9BVTcO01MeRJ3RYdJ3EjLuyomCj7oMI80Wggb16EOLWWAvTx6iJYgIIBAnRPwu1S+bq
q/YnNrDNkGmJW43rV/TlfJ/w3ItMMEQfCcWqFwGgyp+O/dA75yt3G4LDFN9QDL40nI/hy+4r8JTh
9lGZ8PoRQtYyDAKkTGcuczPzJP/JOfzeo7EkJKoSmWMkWTyeaqazP7W/xs23SXW+SJD6M05rLKRG
7r36cAmZTafuoJtLo4cjBzqqHtU6u1nRl2CW4H80u6EIT4F+7YWHBBxFn4B/JC0trvQ5SQuyL29X
kMb8tusxoVaczftkcMtMt8ZWcwarov/APUlqVZ3N+TFVs3IX8EQpv2lITL8LvHXo1LbMaREHe/rv
Fw2FTzQjYyYh8O26oFwk67B7XQ==
`pragma protect end_protected
