// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:32:01 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F4pY2UF+4wS6w8veaCONrlEtMiJr5KepOh3p9YlzZA4fZ11clw2EahBW/McOzubu
g1wv0ecxHk1OgT+7jNQLjJNgePhG+ims0lMyQigkr20b2XfwWFa1ciRbdgBd2E8d
8YhuYur1PnbKahia2/3nPrpiFc1J0wMuIc8OAfoEpzw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7264)
j+7YPGH8JeT29RaCj+RBS0yHwy5tILpdt5i7FZ8Al1aN3TjlOmL1hDde0JhCDvAt
oOVgNfXz32CjvtphI2zHz4WyXUAtXRw6JdZt+tP+Zm0fsazvLW8UXETIkm8K6Dfi
iP1Yo1YuMc7fMdt6vD+ELmjcBHv49pz6wlGNJQ0X8+O2F64wU2EBBCYiCeRvai0q
56djUBJ9ceq+JHxul4nkueTOY5jDeWhyPHAfGwkx4De3S2TlRS2jBOZI7UpAT0LX
6zZKQ/Ec1XThODtllwxTzYjXyBKarvFrig7C9jMSQIFHiGAXgVC5qvzQdHO6kobo
GCuvlVOXIwLInYYIG61DAslmhrgnOOFn5lMxRtK+OeWw30kfsb3VTxT2KnIP5xio
RLM2VgrA8A8AetYBQNFHWrJ1xGJvGyIoQdHfwv3s8zKFCoxvxe1zU/Ez9WHuaKpP
vAoy+NPWohKJKA6ywvbGwC5WPTHc+mQrTtvgPsc6MydAdGDqeXq3vsER2GN5stCI
bgQ15AHFSZ8Pa2MEEAQxU6CTSXktRuKHmEhD7TdUhvhVrE8LwFjOrjsDqWL1CaQB
zphER5L7AhBMWtYJLt6UlB0asibT4VsEoeRp6W9GSAhfNGZyE5vldBfmWRRaTaeR
7vA9czJSGG1HUD8Abd8bGXv0Ut75oNh+rCr6ipu79uAu+unUX6hjdLNPDzcsaXMx
40fsQoTUZ8cNmKShkFlld6w6F1vye8TgmxQR7D+NS5NG9Stdw2L5r1MueKq4Y2Mq
CSsRQKTzgEX9zwSVsiZXbh/Q6fkFN4w/a9pJENrR4+f75eY1oO6H4YB9DSZ0lha5
A+xpywam5wPY2guBmSLlJbqC7APIdsqoxZkfAYa+TWYXW9TYQYA9q/0edWYrrqNO
IAIlQ4qivymSM1kcJ+KrVKZmCqjOxAOoo/B94O/Fzv2G88xudHgUDJuf4IKnOH8A
4Ftv811MeYgm1wmMMGeoSzVtdQVe6hZeZC2/vixJ6NQFII+px9mE17RP3Yx9f6Aj
6J46TZAE8bE+CjDQmQo/i/AKYpx2Jzf1dPNFf4bgOLets39w6eXLbDxkHd/4ai8E
ENKCsTNaUdg/pFfZF4jBtMwUm6IlzZKJvQ0/hkMV+zQlqY5zxolDDUWquo7SefL3
snA74dZHiBXYFmg+4i3xHsXwl+060rTHIiRWno7xShbRi/kEdFsVjxEhoUFwAE9T
2XNBC+gCLtJ0tY3FFJ9DFCy5kSYq1uZa1NsPqxuoY18fWeED48gDt54F945TeWD0
M+V1JRZsI3yd35V5WXTaNsTQjQLihTIlN1I3GKHWUhwUuqtpUzNhgBnVeTeM9my3
lkZb8Eb1jLc8QspuGbPjeiIq3SfK86+Q++C5LJInFTyJJt3Z199Hkzu/MQy4qB1I
RcDdluAjbd095oyaDXJoifsS6RP2vj5sq2nVajdmojf7oVbf2fV5j1MdaLlISTcd
GHmO7y2s5PdwFU9t5v+ZPlkj6YjHHtnUFi68jlSkNAeKFNwRfzHer5hlQoIJtzIc
45iIiMyB4uCyiJLcV/1eQyKTlhPKOqZizhp2rQND7Ywnb3vUDaRr9b0fFTNAHcC1
K30svQY29B2GTMeVCWqmzmpO/5aPsMKYWebVOJClOrAJVvUSGBzemj9GR4JYKl7r
HjZSgH9pbXF62oN9AwUuToZMuDGqeBMHl+YqJIdNvCfD5ZQhjx8nO/ur0R4rw3qL
pjhqbny0c0Jv4y65FnrP1vX/kulhtrKqqSKv3d1eQTU35Y0Ce/UxE/wlMRgbSzh0
0SZZbuAFQuX9FEgLK2Ac/MNHlUJseSkf7FrNeGVQOaUeFcJKX4Jptd6x0R9TuNV6
x+xh6jcJcxZ2GU4IsTEfa05qROarJF3h7Mv1pChL7c10WFELlt2bqotAAGrm42/N
f6PoXxH5zd0An5Y4j4UH47YlDLAosFDjX7caMKNrOfcJllkParuWdxCB5SYK/S60
QayazQWnixzo7O9Aq87GE7hCWuPB9+BD5KSmq/pxQOuS8G53T1nlFpQoV1cuo/t+
wtoxrVzZV/HgsBQ9lwpMbkEVdGMdYAFzFSJQ+YqVUOlh3cqT6GZitSfi4M5b8dJW
GpnVJWR7eq0VLNDV5+ycnxgxrDDeDoPGzEPvwt69HlDlMMh28H1DgmaT5MQDYvDL
G9kzwMuKhkAFjXzF4P6c5gRmp/nT95Yaz2Y/yVTNeQiD98+Yf/4Qo8xwkDFNIn9L
/G9UTsZdmVwkaZjgEdj59oEogELTAbl2T39Yw9c6ct+ICWXjDrbo8ukzrZAkCHug
cUA7veNdDxfnDDCCdH0SzzsOZ209KxP1vO+v3r4Z5pIrI9DrUKdlsDn2g4dt+Pwa
sZ3ITWjjcls3hFfmEXRbVRjfbHM2hhYk4vnl6WFx5GFfOS28AB7zXEgGgxlmyBRb
/dmyM/gdceFXlxRfQLuqeCYuwxlLKAgkMi9WDtZTaw2JGcOny364WcZcBTYiKFVM
h6Ivvo4eCa0+Af6ppPHp3JWfDv+X4HL3/LvVQOoNYljS+gP7li0q5ADGgz4PDa9a
KAeWfGQOvG33Sv6PAdwKfWUD9CQMh7aalEj5BG8L7rWCKzeBvawUi1DKmJqmm9n8
2+7fF3tA17rka46vOrdbw9vRRjc//w7G9ShHSaAc1R96Db8X+9RpabQdcmCQ3iyp
w7JF9leiuxttrgmrPLiqQtryC+2m8RB/fk2Cv0yePBiGKHebnS8GG4rFXSinoFkM
uHAVhpz2Q/vzLymBikXMq71qLOq1P0f4erIiWGehrCpiJTSQym57tNLUx1pTUinw
DQpahNHAHVR+2kzRd497YS5d7SOI2CECboflVqToQooi+y2uKOtdbn2lFBoDVrb1
S1z4KxmuLF+2kMJfHrmHvmyu1ZCptm/1ewDAohZwlL6qXoWfodgJc8oedGmpFMmZ
AYOOSmm+0LSCcA+FV+ByGhLp6gPg6kpQAzBuMr2TeGa342whw8DZF5oCPS93oK2s
yaHrGGjpbAR9K9q9qeo6ST+e64dS/fTCIRMaAOuccBuevS+idlFguGOc1dr1o2yJ
T1m6LMvL3nY8FurfqBZEU6s5x1mc7UdcyASW0uMDqjJaljKljPV2+fPY971qqmgE
7O1JXzqjrMx9YTtWDDPxyX5/h6sHUrvuwzHqcbdcA4hupSlXWfQHFLiToIhXyd+k
X/wBH1t36bGKpfcfHFLcnIuYsbUe3BZvS19BLWBHf13c7J7sCjx5VGAFkpQnFVxE
eDtjgBt8SAePOPfJAtKwFTxKBfS/48djRd3jrWgIB1nUPduIIpgGYUUzSWZh6rcx
MZoARLDbDfelrvtW2V19OyJmdgxPHTpM7u7ZJsrAHux+wkXf4VyVo4wYh6w8MMZf
5/iYR/I0c0Afri8RyaGFGim/6svcU5f+nukjd7B7gG8UqhWlrSnelBVQWjMeE0yB
XZkixORF/u3MsX4OVr+g+BQPW7uqAYZdCHdkrRwP4FmPrTxJjHfPfY5UKD4kSdVz
K0o32hIkkjlpEclbn1D+27Aip3plIWh/YmzB+zSoJ3MLVhjl8hIZAbVwbGyuKyiu
1YjewZ4cqWOj7mPcdqldAU/foVlUM9v6HUPdIjnFWTGI5JrSmrdxzcfkRsDUOJX2
xT29tXvVk0LoI+LOqwK8etzUnwI+sGdwNpkXfZmOiWS8O0u+prVn3buKkPfrM2bB
GyGKGrph3AsH90peYsqIVp3qHiDXg5qOOYlhSm8x+MhDDuCTcuMJrOY/gqX2i/o+
xw9H85fOyTquw184AodsojMe9iD5xsxDgQ5CWJuZxc9l5CADgrZ18bK3XiA45kx0
9kvGCzru25ctrbCMs2YXYcpmPqJPFojDYeYnHVVXi8O0PzOaZgiMee92LFVTHTRu
E1Iu8DBTgbmrFHiBVPdjh5Yr1HHpjHQxaLq/UwBsg7Ql7YjMVE8S0/RsIyMlD/w1
zILOXFoDLni5jOmG1NbD5qyaT4q3qlffveI5cwkOCsvcDFjIGV1Bjn3Z7kzwqNFT
gf7cU9GNG5OUe7OCsJOXhkhpOeh8vhaqDzRiKPin60VG2pyqswULvVw9NLQQumYa
6f0wso15N0jndWv0IGtPS6PkZa4m3RdLBBZkmaA923XIdHGsuZZJWnBNydA4qW7K
77PSaX0c4rdR5GHwSelAgb56czP1R2vLgjuTA8a3E+97+CGNYsQm1y23lOvY0xJd
qaTpX29srvpgSA15CYRUmyMZvUtWQ1j8A+BcvbDposzmVJMat2yRwDS+00OPxS9o
cqeDW+mnyHJXWLCSxBW5HLCvfCSYC2E+56UnNtvZ9+Roi42lfG90cYQrMnZQdP03
3/dVyqD1TWafZ3ePGZ3v+cbj6vfnELn8iIJP15WwMcBi3bd47F+Ramgof0D59Nwu
pHOVNiS2mPRp2/73HNZnkzFFns1MWk4EGAh0ODH5G9DwgQ1nxxmzVR6GcIrz+a8p
rwaeyl7xnB+tTdfIE2lOL2f56a1qD2SchXV7O6qiyTsTeCvP4wWSnA7l5EI6AFQZ
DSln+671Zuglc9+XWV54XV2DthPZds4f74k+jgd5q39NozIShznLV4+UYLf3OTaP
IC3D03zuCwYTQJ46D1neTtrMXXkM6msWFbk4AnM5zDw5GCoAP97aIrNhWxjWsox9
cC5qFUvv0+7+5z82kXHU4ZkN0TyyBM2f40MYmv35zPNc5TSa2bcHqBdg8qYCoDb3
hiS0JJy6QwlBstypSQ0jx+NOhXpx4InGgmkA1c2+dDIz9nKFGxvlFPllrasB+fyV
NWmhoIfJat1OfsgHVF5KAnWScreaQ9EEgQsD+TzeHzNWiy3HduDatSl4PMRtLGma
l1AMakUAMZXqqsr2/M+WmAHr6gim9nVGs6TsUdfr8y3L7z+sJgvc5jRX3VCtPU/1
pXhrzbaeuQnv1/CezxcW0im+X5UfcC3fwH0U/6sQKKMBrj1KpeH8BeiSC+Sx9FI/
e7vynWHKmzckawuLqj6menp2MDxnPplywj6v5Xcd8W8XvbIbU0g91vrQjQBjZmoo
mNUjX3UQBfbenwdhCSrNbueLMKIcSpEaxS0Pn0cvycs00WMvdgsM29894qwZBjbC
VHbSKuLr9943Zt6ffp+PvHwxqEPUQVkDHPSyuwRvMtt95YfzGS+ugGFL+jWBs0yS
K3IpEuPieT72IGoWA4OwhBbu3dzbjOF0QRRaUbMEvuD7MH5NU4702O3Jx4PhVsNc
Ymslik8AxqskuMZ0fbxr+qRgpg5QgMIdcmALA+WdMhC/HTdm9ZEIa6XCPg2vuoBM
gGQqTI/40W20xC5+EtTDaGt7TL+tsISFMmmtVehWP+eHLHSPwkJzLJy+ojxtpXj+
fCG2ItYC3AX6jtlSMbACjPl6pxfdJp3uFFMs5G7PupIPuHU4HpJoPke2LmkAoVNv
NYrpReEcQ7jGEhYhIyzS1gTzovB+k2rPEfsoCQnY50G7DZKNogB7FSUFfdjgZ6fG
QmzPx5ZPbGEgdqOBAdwstJXd0J/DSlX0vFhJeyH2NzDREoEAhSu3tJE+RHAdFWaL
BHkldcsoHgg+cnrPBVlLL54tqI11XfQPdFgd628hGoJCPODFpWDKbCr/yee1WoiI
IpkKaqXfcc3e8c7NgoxtTwyxPATeKk8Qh9VRdH1EpfDEXgNuxBxwzO1Kr+9hT/jD
Huc5gB8J+fPhJvCBJLSwaFXMpKnq55YjRsvg1Osouw4HiPKH3XdgxsGm3SuYXvse
wItdAxCUx1i7IDibpBh4R7li55+FJWOkV9z/Kogn4glfgWD+cW2VxNFaXLs0jf1k
NB7dWzQdyicBkK78Ye+hnEb9m70Kc2XSrtyvGIawKSwPscFNoyjwm3YmFRVRPj+/
X+309RFW7S2zLAQylBYQ9OiCs6RKDZE7M7yzB6sbO4xELlFnvXuoSash0P5PCFyG
hC9E57V9IKkBLyX9c6dOelvE0vz9TxLddPX+5CLjQkT6PR9o94ZzHQ0ZW+PZ4rb1
ANaeZtpFIfj1Beo0tNxiq4KxBHGnas0RiPL7Qx8s9VgNLtcO+isZ6q3gjLGKdqPX
C1+CTH4rRSFn/pyBHijLBxobADs8GPBNS+Idi0++i9OGceupT6ezgpfz52bq8Ya3
PDKXzxbLw8SpjEd0o1xzPWaeeLxcpwiYeVy/acpgpC9tOOfV+ZFDGKHgroBp8N73
HBUDbF/aVjDBmmMretynNaGbEcz4s64Ea04FQh7BptuF3WPxX9ajD9HbAYk27t9C
ES1WphbSxQQALTuDkYlJd//+qTjSDL2f+VIwLKXkXhaI9s7Kd/QxCO8rm/lIfYsa
HLiaADNKed0V5s2EN45xxSpjz45MUqdpnY22tj5lCWtBMpFzHtaRrsG71JvgEPz/
RDkwGfH9KVjemJrzumWkExxRODiVVgohLlPu6HuovBzGKjWbxCGaNfcPwzgZ43F7
hqx2G+FD1unUtDwSnluzqc5jPP2XFxZ/qL74LAzzzGIMY2fNtkSWSo4aEKXe90tj
4YEbBgx36p+RU61lZSGUVPNXC5bTLxeH+HfreNTWBtWPoUkISokFW3hzR5or/kKf
UnGOlyeRSCJYJGzcLBD6qAle65eRB4SLUNxWvzYSwipaxn/fA8T20jLy7OwhhGbj
unytjwVcGCcjdzA28fQypjgMDD0A6tM9R2b0gB26BkLfU16VXrLTmdUd/xiVo2kg
fQ0U7Xxeiru9F6B7z+2M7sMzP4eh1COL22kXaMrDYiTkdc+BIOLb/iJRQzWDP6jQ
CrHYuEi17+JMJR/Ovfv0PMdlY67zzJNbTB7Dt+fopLR/M2SvthR9ZsoyOxdisDOM
BvwnI6Gnk7Kbomk7HTUv5ul9VpGK8MebpnQ/wcKoUgQ8KME0tby1OeT/rQSs/SDB
RmI/o/xRR37IboQL2E8POuJDG1FPVJzw7J3E2yYbapcwp033B/V0ioEUVFkKxrzi
/kbTLc68eCisv21QfWqNwlcVh+Ap70rAQZ+Q8mQcxtKOaZRRu/OimsfNEAZkVNMX
ZLGFGCDQxpyD5RyDf6Ht78JzglmnZlE7Uc595WqIk20DNzNL9CYXun9l0/CXMavr
7btSyYQGs6zwpcImx0pwebdHlL6j3iI8rSxRl0H8ryfDAVKqIHTwwA6Gs67CPV99
0KAkCOsMvy0BFwPG+lKWRmGSJkw5ix/aU+UUXD3fsUnKhJuQQ8GvESLFQhlanH2n
dPzPYTXbZHfN6dPEfwL5Gm6SLcF/UoyZ3C6O0jcyIw3W+irTNcPEL4ZAtbB7lrAS
uw4jwjhWpGOlGUVezf1ofDGgOnTcwqWfTRIwFyoqEbuF4bE5Or34zmNIzVhq5Eao
cYt0wx3NrOEAvewbe0N2Qn/yYcHJgHYVl3lI91jzH8orXeINex4UzW0EBR46W8md
zyaRKw/iuqCEVIrUTpw6EIP/1jxPsuzK/k1CDwmc+SYPc7AEFYYAVh+RmscjcEZn
0Fdu6KPjWUjsEfXO6y6SGtFz4yozZ7+YjzV5jNnVMOZ7VHf2zEaIwC+BbPOePR9g
pHsIdCdPJl0ZIBAiZg62+2oIJg53UJBBmVKV9Ph+hxpXRQ/1+eCYQxMkMfH5KYF6
hgx0wRIFpHhaJ5C3+Nl7Ic13LddWNe3KLoWfxOzEtCYjjMRnYe90h9K9UUZ4aTp5
rF0+b/TH7gVjkJ2y53yeUg5GGnlax9X5edoh3MI+un5Af4t4D+Q+LbdQ/lhlqyEg
5XcVpBk9hJfmDb89GQZaDuFywVpRGz0Hx8hb2ilfb7bywcVS10U9TVNoO3ETA5u0
E/Nv+Yq6hUWGpCFaDP6qtBJt5KX22qNKWzUYVKVu78cMZwsqApKks75IQVApCaPh
MGTDlFDSQzkLd/m/ZevCeyo0bVEFQvZUwZ+rNHBAfK0FZkZ64d4QFwcjNhxU+G1x
eVcR6em1eeIqfFhNldK4Ifetg+jDhI5aRiddGS0m4yEjS3DkQ8NSDpFgnjRj/7y7
CgrKyG81IBq+Fc9tZbSseQOGakGvlHbeAheNuHeLIA04v7O+Kh6oVvtZpBvHbg3L
triAL5mIB1kGFdJ/kioNY37NvpkiM7ePms4QpQmGQ9eCiS/Mq9EznLux9Tn4X9t7
YW8FIbFcxgOB7XTqvapL/w8/c9h1Df4vp5vtt/zyQWWIUhzcE6JroE+gGXrl0kiV
GQL0EX7/QFsSexXJ0vV0A3j3F8hnbwX58omw+TyENOIO+VwyhN4+B7njkhnagNL9
ZGES16lMwwRnaDGlxhL/8EsNvo8VoMcZ/6vvq6lcD2HdHi92hAW+evM+ZS38lNDN
RM38o1oYez8CN5u8my7XGL5pjMnuwkKK97kqN6WWnEjbxgeLegFZoau+AaBOD7zK
Y+dlxGoe1v42EtxzLTQNFD0Ej2iQLNI0H/KAlAHqsPsKH/Die99FOefguw96BZBj
gxqrrIGrI1shGmCTyEvuBbbJd1dlq6DmlW3/7RnWtxSXxDRVkq7J07Yr/oAGSW8Y
ckwfbbxyCBJPzIVod1k4I9VZNaQwn85/1oJL3mmfllUgJVDtsK1tT7xHs6/ZqsFs
+WY9rTsHu2Y43bW+2zsvi3BQT6HE887W4YU3Rx3XrrpIS89e2PTaXGuy+YfH/EoI
t4b61H8xE8xw3/js/YOT7uO+YDlsBbFuTBdR8bot8PGOaPdMbuTPYB4Nt3OdqZYp
F03o4YV2bsr8kmmZW9eL1lanx1FPhn5vCi3mFVfejysq4Do/WUSONZEuQXVHs31i
4cVMrCtT03ZvtJgaygShct7F87QTAFp8gqcln0SvnJfG8fcutp+aftJDR6jbh++F
pLovbMGGgxRYH4uR9AApPmPEhS+w7obDnnT6qruqc2a1ebYAs/Sw78jnvjX8KWRY
7BsoHFIXocxynFnLDWLVwiehzJpMSJUXwSsjZgMlQ6raKry6Ak64QP+QZPJW41AE
tG1HwhiNLbqH+FX0IuhsmJFfQUZLAjCXb/Fd6FS3RYEfkUUT51wPqx+yf4pWvKtc
w1fkKtD+9UgkVipWDZaTtyvAuK8tzHEX7CTTJxpvMBdM6wcdrWOE/k6qdpOb4dul
dmAbAB4OUEAoX/sFUd7Sn6a0rwG01mTRXnJBC1HuhY/0LVftVvW7H31KH/ASmN1W
hBLJPE6u8giDnhLrwp5ukcYIAE6dTKlc3hcCs8g9h9eHHyEXLHcw+ei9JoH8+5gl
QuKTGIZl/+vN/6PmtVfP8Kx3D1TbErH95LEF84w/kR1JTtguFpZvfLYoSkxkdhqT
3OsQFLnMFwAM0QDMwA/UGOsPeSo4c2fGqpsQfIRKamD1OsbTbv2Z0xVs5mU0Wcjn
HWPK4csHQRf6vpYbsc3aYvog7IDots5BuR3c9Mes99LL3BZxKjFqwoR4B/vDMzWX
0QDqwqjjilFFtu+Eu9XNTbbMsS4SpOQs37kYOPyRchTyKgmrLA20oASYJRrdo3y3
0V7NXqoqHcwsLe/WNNI+2XTT3aCOQjXJ34j4yB7swxybqllGTDtMRz4KAq04BxWk
nir2QZv0A2Eb3/+hUtY/mzD2398YGECbfYbDCtitTHz2+P5eUa1LV39v5f/NJwbo
P2ABBpDCBoR6phMa4RcLOstYNQC1QOV90+cy5V4sHahn/4HuMcLI3c78/K4cHWd2
Cn3KDQQ2hSHpPFm+Hm3o4A==
`pragma protect end_protected
