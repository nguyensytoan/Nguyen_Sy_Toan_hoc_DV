// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:32:02 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Rnirmn7l42uZcWVcWRhnI+0bmg7trRrZAPscZqcvzJ/lpz9mZ7RQ+pf0RFbcw4GR
24bnv2o5HhKOCYRxfrRR+58B0QzRw6nrbuWRzhPYaKHCe6I2GcfVYMngVZ2JT8Z1
h6tBm32v8RyhS35r+Wx7S97SeVWmuD96GrZojuW2AdU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13824)
wwFev1EeX6NnpRu7I5c4pp/VofVshcsN/SBCEZw+U+6pKrDNdyOsyIrAilsYGiae
w/fws8fJc1rItU0pucl6j+jMhOlBWpYC0JWGVS4yVzF4n7IUietgYh2pLg1lB6//
WWdgTJV4xUyUSZJuS6nQ2Npe/8MJXytyNmoWtILQcOlrC1Qv0jfdgCGrc/Y4Intt
jMUQGqPAi6EMpvTUgoQP/MWda+i5MXoPBJYb2DGElidv+KScFTbS/434lDeKuAGh
Awti9AHmHIwPumQQvXmRWE37A1BloFwsBEmcYAKDsjZKsw8pjrl39U0XRLo1wHPG
ln/cpzA18c/Gpb/WdpD0cKl8by15GGS0xutpGXbo/H3iL00CZ/SR7N/gR676ECTp
1d8Llq2sZ8ssSvpMRrPy6cAqEaF8j1NFWB4xsanVKq43Hf+GMElePgB2gBq90EOa
D4vsmam1Iq8lDzyrhCDtaeUXhbq8EF0xwt69c4uI7FPnh45HQUak1O2fM5Hs1vI1
HB5yDEfv/V0ffMWwufG3yf6Y7tUK0X7ogtr6YgVj0agy+DFCALeyV1eZcscs2J5r
VyPTGEF+SRERcK1znrZfIXtPZt5a25bCQFl9md8jE0S22mIwbW0yrpssQBgTkvhV
9TzZVQORviAuXq/zTpQ22HkL9Jf1T5Ech+X9Mt6+mCwmPCafjlsKCeHCk1Cd6rHb
R8RkCuRJtkZE1XbYAfANetBWGpnNqKbS5fpxL/+SRi5UrrrlPoVgLM9trflrHi4K
oV+ntSws5Y7rG4UPx3OneS8oTXkCtHXsaw/+Z3x2O+VX4uAcR7BJK84mlLgl0tVi
pMCVLZ9XoBFeYNiimXkkXAPZe+2dsvdc90tlm8ICp1S+NdSoPYOn4GDCWxX/Eucq
H4P96U+irJWjict31YFHXJ+2RPH6bR3Cc08xhhsdDBGesl/f3EyOW4Kkinhio/ng
4roktRNl0Teoxlw2PSN5MKsDGAJM/y6lvJcK6W2+g33GE8gu2bXQF2cp5auFgX9N
KaZrEoaE2e5qEZe1n7vpjVXqqgPI++yhE/xlyMZniWgAHYArmHsYxRFq5A1zZq/9
Dji/YOonJH68I5rx9E56/PpQw0TY04CkT+WH1KvkiFVHfgXhbKYzZWcpa0Bq/M/Y
5JwU49vfyeZJWsAjPcbAGXS9VPxz+44534hbUTpOmBTIMLRL/hpKPDoQGijw7ZCh
t5dlk68KcWL7Psy6PBYENmfrqE5z8+HKVh42ixocXo9NHfPmPlHddwPMkqe++Pke
76sDjHQuW++fyiC1OT5zJ8GasJDFPIqg/ZYelTRcVfUhfkQ68O8M0nP0s0hlRTT1
caED+IS7uUm2rUmhqseJ+Ik6CUvaF3myy7+G6KYDeJneiI1DcJuoAuwNBCeVXQoj
+8u09x0WBiyz0hW/1R8RMaKKxczPSS9sN7SaQjJye16Yb37ynXdmxOxzQzvd6n04
b+JZQzOp6qQIZu4HePPRsxALRHI344kZOO8YYRg1Dyr++YDgft6GKasD7iu3jZUF
o+/9t2e0nk1gmJVCqzaX161Heax7l4lhaN335+DKlxPFm1FLqZcaE0J5cb5K86+S
Ywkt/0guuhPLw68swHZnZ7LtRo+bQi2yz7XqLyjt2bYYvNjx280DN3L7tBeJj0T2
xkzU8FbXVpBMscasIg81rIeCuSb3tVJw4NcRf4Q0JJA28/4JxUGBbdlYv33b1u8O
PDQRrOtQitnHIyx8CMwu4DC/1eFoiVBB6/29gNf5jnuvTIeHxb5sexKRzQHSJwca
UCkNuPslC0+MsDoWo63RxO1zoMBoG0KUB5fLWVmzcFc6+xiBgZlxddEROrzYQbDc
Zbh6B8MwwIh7jgxQkOKB45WFIh+1q54N2Qzr+z2ZGCHvQrJGIZN/UAWiEryx0z4X
D3mK5UOh5ae7VfVHQblBGGYekGTqezqMw4y45u9r1a/H/sSBXMesmT01UXzc3T8l
GtmkifMlEMtl7mr+ftzAYvt3NxRC4j7CIWeNVf1/l2V9WZg+BAzfDjykTli1FxoW
SRQxcH4bqR+Xq9Ppjv162ZTLZjsxIBACnhUI/fvBqD2rqLt688Me2XDeEYhuFfiR
06B+2Yk+dHi95suPSJQN1UtYYX9cmWWHVwABXn++U6OW2x2tPzNV/CvjEVVt8Zq9
nFBey6xlY8gramQ6Zyf7AXJowzNlgCWyHNW2NO0o3eSojy56m922XqjB1s46/2Jo
LrTT0Q3IwvKIzuq9JgLl8WjSgXxM+uau3w9/2CPWomaC7VXUWGK96BBjdDe6KT1M
IIT/O2Ejl97SXsP8oodRQO7N8A0uwuNg6j2hKPIlOtZL9dKWJysYb/tN2nUJmRLZ
BrMtblDSGtZctpeXnc8BLIt70ViV79TAbODcZ9n/tym6DDJtsIAS5vNSPeWo5DCC
hbqkWyDcdsJqeKPY9ZGh659y2XI1regV0lcVuc9hiL5UR2qROOa2JGvOZQbZ/nOP
GI2B4xH1bC2obf61zJI1tgOf8gWZEvL/CFNyuwKRGEBbT8oPM5SFX0eTjDUvQaJ2
H5t4VK3roSLiNauIRTUPUt0uESnaIPi8ZX4Za0b10tofjBkL28oqWtgtgK/me35/
HpnhOUcZCgqsIeCVmamdvC9JGdv3UwDRBqXTFEkTl4S1RGJeW/jlTt0Qix7HYCRU
/co0RbBfKb2N6eu/ACeXSJRCC8BmeY68X0JNkvHBE72vyuxrlHw3C+2Rv3ktIVON
HQgRl4R5xg1IX+G0lWXo1vtPQ3jLY4+G5p5XfvVAS1KYaShOCJnrDSyvCJDCz05a
QMehAA1Ed0eW/8oVb3sA2UURvvgKe6GPLp7IA/GxFojIgY1cd/ohvKrTqjyuHEoI
KBatFk4OTGJ4kbrF7M68Dveis8ckoH8sYEDrrMnjn5bIHZN46GXlBk5iYj9WjU0N
qhCZviikJ+sViVZxw+2m43ZYYqFpl+d5YSY6I7hKoA+dYWHL6OgBTN2W5iERUK5C
eB/uW0zL7jNB16gr67PhFaEN+DOmSjvXOadcGIIbc5c0wVwrNTJwU9h2KNhQfGg1
41E3oLZSJrvWmBYfFrOLV7RYK+LHwqp+08SDpJ8dtqRGxEVNC/0Fth1e2N7IQNl/
HCBkrrhINa+81Yy8EsJWPoNIk42KtOynVS3WQr9ynBg9yGmDFVTo+A7PhvxY53ym
JG+d2iJJ+vbcj27SZhJzUf+FKxEmN4c6AfzRagLZuW0Hu9LNOnshM3DzKIz1LLOR
jT51ypfsuNTRok10fyFV4OdUVIBSrlbn2ZhsHk3wc74B990xYQTOMEqNwXJb+hwP
0lDkX7XHRSS2KZyZk8apXScvnNUhpWpackQSv93hyvAANtZPYcev0DVMEtwyUfk7
JDz5uNvaGXNJh8TXgfOcBDPXQs4quqVj7QP2dNZ6Joel0rjk+MTJQx4MDFtny4+8
Lyfprncw0BHy6B1sFgIPbQS3IMB3jdm2uwK8m5NrJwodN6JT7yvs44f+SUxjSfSr
oW/aEin97JvZsbyYmTHGOUQtPGlkNkJxDDOwBGwBX7eomLSCm8BDdJYw2Z3kA1+z
PNQryIAyxUn4OfiKtzvpeKAZuJpxn9KltCGfIs+EOVkeZR+LK7VrnGrdlGYqqeYM
YypJOu6RWus8lwn+NXV+Be+/ymjliDONPVmi4EG/pnTY/C1OyLpnfSuZ5GFF8ekF
heRG/hpBBlLMjp9kyfskHE1vPUBsicWW9EesJEOgACSJjtNa0gVvrtY+QDfFqoZY
tnyravk/j4fXpFPNfDJvvRdjfDMvIEJUmDYKJTZw1JYUqtwlC98yGewJ8IaBKA27
3GJhn7LqgZvo4JeArv+IuthQ3V2Chb7fk5YZbIPR7P2auS9H9op7/Azg7HY1eWqg
OAhiM1e6WPak0Md0ML1qDCjZ2xmVTtMCf1Cgxi6B/sAJCkSujruTlrYy6OoBsEhh
KHUcso77BBY/Ivz3j+Ba4nQV1cYsBv8J4/OyedTkCGYTSoqyswXc57UKaMrNnU2d
3KFs/lV4Hx06XVjtIMY3lWFfGsqII++wGoA0DbAUVB1dA+a2RcZ/6lEtXjTVvQio
ZZ4uO8y83J/eyWggrv87FmfrZx9p+LXc+PLHY34YbZYmocqok6qbptYRxcBu+YGJ
scxpGhsYwsaM0Qx49AZI1m7mwSGKL9tndrNbqHQY5Ye0qmFJZw7nRJ4yVj2gECJX
cuq6zEw+1FkKO3SWOW/xv0Tntz1CnoQRCGKbKJSwzS8cY7ee4yE2SgkYWz1Z55DX
orLtV36V3p49QFtLMkPM8rCMzcz4dqDnjb1QZiX8834Wka4UQatinun3IZ8Ly468
wx4tMOyB4DoE4XEFF/sza6vnVXqCB8TZVzxM4+68vyx/ebyMvGPwtLQyw13e7z46
9onymndrVFsw1FLwUnVljaukEzvLROZne1fh/rNa05nez7HzVmrRM/bgJZbHMu4s
ltxMSlyL2MDXWvw19cyq0mjaElpjIoleW1uuGZ5VQwjh9Cb1O6aTY8uqbFwMzrZ/
06Q9/B1iKVuBnghQmR8yUIXSCN1+Bp236WINAAHoRPsQuTUMQ4MmQe5He8qkZ/ZX
h6CbrQojwy6a8Dqk4yvfVIR35MkCCM+OBN8ieFYCQDfeX6lugLqWAD1wMz4UFUJi
XM6IszBBJT8ZnCWV/TKNgLLwCMZyfcyrUlHSYDeFzh6nBO45HOZOYTml2cRxxMZu
pFNlP697oRYmP2I7R/cSvprDYBJY89tyFs+4tqhNkd5NmraAM5Ua+pReFERinpuz
sCOwq4Jn6XKFpRPHkVq3GvZbNOMiM0lleIA1rsCDVpZRjmvXfry5rkFgRZKtznW7
m03bf1aqGDNtn/dlOjc/IkTj5q/I07RJY4cfwtd0Jz5GKIVpjJcmes8rTVL40DjC
FNpRDF2xpTjXNqF/ywQqpHkahcMrg3Z7EOesH/r8R+9w1/HPXfmxReLyGigIQHWX
KvbT0OQqIODCZDt68L86+jWLVSJAt8BHvxxfZnH46p2SbEQwO5VOBuBV/RvukV22
/XCqT9eh8vWh7mIBCx96QklzrENwoEywFF8xs8zOnxGzkuAHycq2LzDtDhJHD4B3
fcnJKwxY6Z74b7bQizq4oV00C9FZsjB0GHOHtrK7WdsMNdWl1pjdpGUkJOYPVZm3
EwYgMUa2WTyu4haANJhTFUnV/xxEN/b/Um2Cj0NDwxlvC/Cx2vZ14BD1fBi8wBdn
ue242Yr4kzPqAb8dSrqCKpI0wCbSIs4F3Cjqov1gAJ+DnRL3FgwqpxdSsesjuEbv
F+77uASW+qni4moZbUi68TYFtgVhrHnQlIXmQ3XX/t4TnfcN/tD7fEt9Pikwq6U8
ngzafKzxRJrCo+pvPwAVYbMh10vJdiqVdCuYwfAdpL8uYQhHy3cGlDod4/Pm3blm
Sb4TqG3PVU2MFlT0dtJD+gLrI29nXaCqKeIT3vyBTSOIL6iURiUA5lrlER0zp0xH
C/Sn/RhwUAysOEpJKUWln9klCf/zJwDa7Dr6klUARKAgDxDfC6MagYxuHRLWP60j
PPEx1X0pfhsQcv6ksU1FslH2Jc1GyUTKhr44t/U1bBPitfv/Q9zlW6ql/C+9PUx0
EswABojcQ+6W9uDXgu966unhmqOerdZiJoSajlNafQ86oLU6bmViJ0yXbz1W53d/
xsyoKIrYldTmoCeoHtAcEqGL6usSs711jwcwBCmAsKHXw40p5jKtLT9C2kdmOEYR
DOcsufBLY3IYJf7zPzj7gXG95phbmL81+AAms6E4mgi+Nzn5oraEAwcdb/L1A7Fp
5R6pQgc1XFld9MhlKFPwd2uu1xBhH+jCGoJXjOwli9J3X24dhTTlRYGaEpkl2BzI
Hxvo8lmFyFo98zBwGNVMph6A22FXAnoEs/UXjSN9RR4PBDS57YvbUBzg8+yvNc2y
weCEE8KH3EfmQ+tiFucvG7fb7FG09Vja2GvhQYNv+2bChP47WyehWNiy8wEl/g25
O4Fezw077djHIDa5+roG/myHbtlsb2SIY0JB7WsxeOgdSAnDUfqxzj72mYsArNZZ
Di825UR7Km2EqhBT1shNLci0woIUSfcHS0saPURBT6RudwJow7N3mRUC7lvcE7hQ
sI6H4czr5hhNpk5pzcEy//zI5XKmEPRqcbwQFktGAwwQ3Q2W71bj4qtpNJA1tuwL
Aa4mmNoId2psYtsJlXBDXdotHqDkXbS1Re6gGqoT/YFWwGx4rCpzyexf4otkU5zY
D2lVqb8ANYdJb/sdB7yrC49BWJfGZVlqDdaUf/Wu0wzIupeud/GCZQej2sFwthgR
O8KQ2IKxYWiaNGXR+ZhayLv8BU7vfQlohdQ+nRvAegEWzMoDXXnd6zync5Fcq0ym
LkCUuQ8Koi2RamEr1JWj+sMb0z7vyKUX99KmlFL8HUjtvi6M6yVNEe5xub66TuWC
ogHHOCn9qbRbb4SO9zKCPGSQDNYHLpjMy+97qnHkatp7JTbLtcMpmPNOdetUWOhK
e3hkoaJ8Hx8ao44hvH6dvFXpbhvnCKx0j/tmQxMK5OpYQXEYMnd6lzmaZj63ywNf
IIMkWu/ract9Vg3LJMt01Z7FUv0LB+sVW3Lk7rZ7yK5EXJMvEsMkJ8Fkn7Ju1hxQ
T3YmTD/m1xciYx3QH0qr656QixspCW2dDoE4gfADb7WmyjhDNty/7ZV/rOYUsv6M
ha7/9DOnZ6zkaj03cAQpkftMZoi57odx2clfhqwYBh089Pp1314NJnEg1MeNvgGj
S6u79rdvqNnXtsz48e9BWd33XLdAKHWabnGUu1nF2dOW160mx9PqMVCVcqssgjrQ
oC1FCK5m/5deyB+BXqagZADOGnxNGql+Iy8ze4Sj79awL463fX2KmZcQ6shlSxOd
59aOY1RvHMfCao5JOgfo2m9/HrDdQ6zfc38N4SBin/5C/uECVYUn1aVhPEgjDJgY
5eS+WhEXQdU586JjW6IPd+NupJ248Y7xKNPXh2Z1C6CFkrK6NDTej7o7L5zdwAfd
GZUJh/eCMp3FPd3ioZI9ruQSmeXACoFhNy/di4I7ngVPsXhqaeyiUPa6TqiGpd3g
sOd5SVBeOOczkMH2iYDe1C+s48XQ7HsLR0AQAMwYlB9XS0soFYlx3MWmjpzFeESh
Q6Yh08K3ZjylQP+mgbocO/xRyrT1SBnxqu3xQtY2Ncv9axubYG8fZH4VwB5KHNAd
Eh6UrDO2/DlB5h9zHjyI+P1DsbVVWp0Ut2XIMWil0gTCt8BzyI2wAq0CV20i8S81
rM2Hc06dd3VIkqnmMXJLwRMlJtU/lrVZZe3hYTRWCC8xxkRFV8l1/Iq/z3sbvNZF
4MOHogzRKAmYzsbFha0oFbv2YICFuLo+3ua2JQAAt6aVtesXHGGcqIQ+F9EBU2md
WKYoLNw6MOWIP6hyiQke048yuypd/kMnDNgzgI1MNKiHjN3UppeES6XkEWejvIt7
1AO3QdqrKcJKn1Focd7N0OtiIZRlw7YuHDRqaYy+Q7Fbgu3ymtxAj/QGmlkwF25f
97cGdZgzk+pKhC5jIPjcwCgfCCnU1rBaEpPFwhK/F5PR29Ur2V29qTZN1r9L3FcJ
XvQuStv7Ed2aYOmKK+DyjUe0KbHplPFj5MkruFGkU5qYUZoeCfV9jtKbIel3+oEP
HLMly1vod1iHvBqEivufHzSZDTcQh2tfwR5si/NchH3kV9kkCSjOmcx6KShmC2u+
dC5fAl7nTUPHFFR+TPHvuZ1tdfqkjfATeQnlBlOJxQZRETx5WDebTj9SS1Ibklth
xYB4fsUpYiIP/JONHm/D28NAnm5+10NruSxd3O0HN9p5+FSiYWYIMU/WUYEWhNGc
JoC/4uU5Ye8oKgBBx2RfYPY5DZi+V/ef8mwIqE2AwfWMf9ev+rWedoXdVpc4g7Ex
xItyak43TQQR4J/YnJKLHHIcE1DZm1YeIqV1yvCAtO0KOP+NRUGDDkfla00Jc34I
1PSKZ9xGXja2sI+VoGnp0oDi3l1vksyi3puP4XG/LZEtH/0fpY2j3vCQhfofwJJy
q6/SBZA46Bd0r4LRPFBMfkfvpsRt9UHq4RUxwanHs8A3c6lBhI0RUh84Rn+eaNLQ
iDeATDjZ2DyT1ipSzNQ0iwDbOF8TA2BBzMH1yhuaLow51WkwnZQwte/lXIcG2ykv
yLf/jLXPiGjNA0az/HdkXqq2hsOOox6QrU0PsvE78CvnJyiPyhVFi5F3ShTPvCBB
Vx7Tzpdp+gJ62/5RWG/4ZS5eTzOp3UrKMCRASbCnSQnNtaU1dKGw5ZDzu0DF0DnE
gdemawRIxOnr2cinHukMX/umNOtML1ajYt2lZBKuK8BJPBr6RdAPtvsf0NBjvXyx
Otm2P/VbAay/KTY8flrFtqkGF6ETb3QDrOuX5GlvvEwm1+vXmyyyxm+6we1K5kxj
kLISfsnxT2mukg7diqYYaS2+D4AjQWbJs+gDHJxRhTekVkV/XUCq6qTorKbiKgas
0BMveuWhkVl9Uf4Sq74RNHFPn65I4ISpiINuySAaTRrOIDInIWqPKmUQpyo+rmUF
Jm+OiWgyso5+T6SbU44NLAWZe+u6hZC/v85cM3pi2MMu0DRJk9ikQqJhcJ+MGSjx
w6eEAzIafLKzN2TeHMhjKfyThZg19w4lJE1IrL69Kpfjj9PjcmtZ9REnwcw392OH
e1MvAOoOnkJGBU3hlbbOez6VJuHwQ5o81WIlNdBl6+JS2QjLSrTqBIrCrjqIKguq
1IO/RBhoV+Gtm/72XLf5zf7eja7DvIHwRdUTeRHxtMgVUAlKbQgpO1ivJDldDuKm
Hk+BCUs0/matZGWWN3xurpqZg+79vnd0iMk8gLZ4fqRWqkfTIiHB94RJcnN4iLg6
XdMpTjG3ctoJluEXKZUiqXo4tUFv/yc4CNWGnR1P7lZj8ejFWw7fS/lqirdkLmpG
U8gzv1McTDn6hXoiim4impf9gN5EtYil5Jgwdr4eS2HCR+DyugPNaBRaBl10yJYZ
UNPVS9cBIgTuxSCYMZ0xGGYjPhI0tGj63zE6CmhEaprpgOIxPRtJRLN9XLTN+lb3
uYWLwWXbRw1jR6kpMVwGzSSEx46TLjkL+sc2EG7Lz+6irh3pFKyyunrL0u85G5+b
DeObqQxUr/pdmUu5Bpv8w3KW/pub9vZuXLaUQoFOYkrc0xHkuEfgZz84OnyyPqGT
m5oF+vCAiJKo584oXqMsB9a4WG9ALbN3C/kFgq5B+ZmZOL3JC4txHe1M8fLpexLH
68lrJohWR9nc7F6Krs4z/yVwVd4HzmNeHWnCS/N3c6Kxn0hnLyPaGMomW9Q1VEtO
tM4+t34wg5TgMajeDFv/+MzTK9hWdOxEMp3DP8QIqrRkuOs5iVoO9h4OZUPTWzr+
DdpR1nnvBO2+/HuTBBqhQi4OTaz1hIm/IvNilXmUK+YqejoFyVtrra9Om/dBjN5P
Za6l5Uz20D+dxdEO3m2z2vlpTv6ip3EqUU+U2uTnnPP6FNdzFYOhbtoEA4NVPVFI
mxFAkT6nw3Fly+G20kD5C6Tlh3za5vzDxBVFGFGr82c7VriuFsCGKjbZLaLulhkv
jvZVwXxhDVMmBeGPMQOSgoHxEjw/AkKrWp2/5e2bGRujGAOEBv1LJAoqHEZQsqS+
RZi12qgLffS7F0dfa8P+uEY8oUxJhXelaa+7sZUprIdXXvUndzXHabwujUBF/sJ4
k1H9QeLDzu4byNg/Sn551TlYZy61Wy7ua6vTt8aSFpKtrJJQcNnw6Jf4QOokfVox
hkXWR1k6XLIj/BsfgA5swLfsbx0hNMWHbHuJGruAxeuO8G3Hv/SaBQLuDnSAFRgv
5IWJ9gLvrbDGIl7fimoeu//CARD+62jB5fQXnnPIn4BFJuqBVf3ZPH1S/za8IMfx
YZugtoy9slVpzoN7/kGUyR2Y0CuxgBBmAfczu+BgXC7rSpAoG940TtG+TF1ecun7
OFxBOCQeSsQvXmI5W13C73llMYs3xLiaVhwBJOyKF7vTreMKeI5kK9vIceZqK2TI
yjdVjho18/fkxoUF0NJaraw5VQw7kToTx+MDsmusC6cdhHNeAi3a24QYXiMTB2Pa
lqRFJ8Hr+ie9nQl/NWUoenqavGq1JHEnK31msey+26bNpWbqMsxfIBawG1wuOeQw
f99/vQDZPDRPjgoMptu0nk0RR8qBJ4Y2SQ8BqcUsmitUhcY6abMaPPm8eQ3aDZgd
YwHav+OljaglGas/coFkQo5WmvL6JYKRK4jmKrFl9sB2Ewu0Bej+uv2aKdrTkkRq
ebKfBC4JP1dQ3wDd4lqbL5N524KcxYfk5ourMmZfND5/Ptxijfk/S0RWtaPRXBHm
CLYxWLGu64mQK7PCYwfEJbV2YoKVahF4BiY17J4cHnoQmHtf8R8JKD6C8sdi8Q8f
GdYyuj5HE2VERUbwJO+j4NMC048itcEdYNXGJEurl5aPsx0flFXE4zTpYxTJZ4KH
ahApL8z6wKNhJjonTmMePH8Gi6Ts3IVwgg05yvfSOYC4HE61dVMiP31mppxRx69M
yU87yL3EHv0VUNzOnLgS4376PuddBYzjdPCdtZFsyiHpC+5+bqukwj6fVWRyOROL
IJA03JFgFJMub48jXNd4C1utAtYrJ7HbZdVynhJ7o2cconm/qCIeiqgRjV2AhzGc
dLyTAmnO65wJSrT6fNauEODtENgkYlXpa/xYbOnuxfJQw/aG/5la9bmX8YWNRl+P
AXpQld9zq/a+S6zKnpPRCK8c0tnP6pKyE5xlz7PCYYPSLkKQjGCUR5GDVHqeVJur
+oONed8uh3VjyIQzQAEHaFX8d6HZxUTufHJiI5U8+TN0iX0gbxqQAOBVhi70F5e5
GFz6eUFlhP6iEH/6ApRmgk+YeQFagY1tXplASBrEqcO4mb6pJUB0DNvcRwh7pE2m
SUX97KCFcle87eNBBol3zMcLR8Hrpc52wm8/JyhzTM5Lexzr7pU6tCXNzTA7Lnp5
ZH3Cq4dYg9DP1MFoR3VrZKL5KFjGUUt+WVDicXCszmxRpZCkwPJQBRgBoTR+UVrz
QnRBRJtwaF2FOfuWdVAFj6/wdIIjif+gtJW7he+teSybtaVo5vutH91dm2phJiG1
dkzaFQMdSRPB4q6CmMsvWmQgHFUWOv9Din1+f7jUXK2pEZeuWL2Lr59efClxDjPM
JWdf9ZaHEWejBX76SyQNSYkJMgRpCE9QW6xWst9as6QyoRCKo+DYJU++B6T8Stob
B17jVGMTNtzpQ6xldRlVCLirNFjCNE8Y4IY56tJCuOK0NAsyBPDKGQ43NANbITQd
JIffVgmPn03Ssnp0T2tlBgnrsrWQ79KrJz8bGt2rOKNhARrfZqOXdIemLaA8DKg5
m6BcEKnefxe5nXSMxGpG44Wfup0je0wbGXuNECBADe85zBK9RFUPjIK17nkzl2H5
OkA+cLJzIiTfAlsVejmZddd+cl4TBp/T4HLDYxwutyw7AIp3d+Dc+z06AOAvaXr5
5I4g++fceaz8ZDy/pXKe/jsw2Mz6RD7mNDIzqmkXov1j1UWQhCbkoJfjgc37CNcB
3oUhxjA1F4/MDLK+I4NwKvkgcZxUwsnlitmL1UkZRRnkTLvEzcGOlcg53386joxT
l0DcNNEPBRPyxCnDN0OZl6DDzd9kSUAkARAgmYHhH1RMdvCIbLsicXWht3PUR7NX
VVLCeQ7d8A2qb22ql80JVKrQ6ZP8K3nohlJWzDq8w5IDp3eBOabgdbJDk702QgKF
PrkAkodDTONZnTIJfdh2bOTUdDg9cLipuJAr5CJo/dkEc5frA8y8WoFJdKTtHL2z
aiMAdV4ud5URF7Xq1sH9+zIUowBPQGUnQMT4fXlNk5T6xPcDS3FJnPr6UQ6LEDaM
UCoAt7RaXXs/Rz01VwZesIZHDXniAJ/llJrLBhJvaHUBz+UM14oCXYNyHEG6xa9k
Sao+4qP+DC2KJH0Ud2eaTWK2xSIQ83y7I4+gh6iKXzOPu40M8IUtJ8F5jSFAd/Qr
lLvxwyD9biQIDdooX+NGzaLO8LNn358EUtj4PX2m56ESodguihNI63bF/gIBIiPr
OzB132ieL/KjYkrm/ATAE2TEeoirNiM2L5lRnmJ95D5G3/6XXFql5mBRUOUfuu1b
ZBNGgrP9eUvt2KiNwh/wqZgh5pWGucO3yrp15aItOaAWQkmsSPXduK5HMF0W7xxD
KgYrSPHNTzhlqAzDVGSH4sof/hfHIfbIxO8UNL99aKUXlPFCi90tCv1ZIf2o8Knt
CudNlz1Lnw/2iuqJYPtNGdX56YzTjUB5ZDOcE1/r0o0RPxN4V2FtLqEl3NLIqf4X
Ty2HxdJJgU/uZ7Mjq5Ls2pFDHOs5U5s/ByQdhs0JNSDHG6WmaaK8EqZX4vzp0BjT
r78pMgDRExciNO4EtqWSPxzTA7X4EWqa6fS24/qZfMg/KWo9NzSOywB98FfuTyb6
gjr8yLlLWrrR61RFaZ3iaW9NltHu9+nfc27Gz+E5eQNQ3117OWrZXkZdf7hzuZMX
aStMhbRF/IhjQgpYqOTSbJsh0GjBceQf2aMHn86i69Wo301C2cwPL2naF1csMLKW
ci21uoMe6/xCDzNtvmVwFwBym99vzSw8cwsGSO3skbPA7r7isTu07jksLX1QNz3l
ozXha6/o41gfTJ1U0W0Aakm2Cs0uUD0CHRn2O4r3FTUbSK2sg0ydJ2awsxms5ffc
BzoEbJOJAHhSmiNFatD0SeH0G3LaOUAZXYk+0sl+64ezPVbl3E5vPgdMjQ1CWBa7
KFpXv9es10jtcTwmw4KJZKHOFlrGEwsndo6dC7wLphR9KpEuiTArX8oBbdvNgnxA
fot7R/4BeVnsDUyS1VR1JBstUvl5J/Bc+QqnZCfmr0x0BXcTlNA8s02kjAZRFenR
roj/g9FG/h8OqxcZh6Muw/je9q2legddy9GFLKOtrQM0b3U6AvY1TwYDVs3uqZKi
COeCMhRAFBJ+lInE4+4FAm7yE63OsIDAs4N4V7esxr7rxNMjMsmzrKeJJH1mVt23
dBPTd89elIfI5/gUOiALledGk1qTIKYDM2DxacVNX+Pze8UVKhmRcq5xcMcYVyN0
/7Wa+zU4kXA4k0zzx/wTWb11y4GyOF43Id0YVIBqPTKiB0aKZlpakZnVsBeki8LK
gnXnMsli2rrlkEn3/9YoOreKniIE8d+ScorXUpZtF/N8pygRDGWJvP7NQn+RLmLk
1+F30xe0ezJ8BOwddXQBqQzkZcqQX7Lq5UEp7FZ5y8cckJXfcIVeN/3u7cC4MbT8
YBI34OzNIDA4KcDGliKLfMhhCJ35IfrnGydkP0eWx0kYCkHukCeHwUAG0B1EunSQ
rhY9dKqpGbZZXqKTGDUk35SoVHxFICcOaWnFuSeLCnHSx5lvwJX9ViM3cCQpGIgd
IbnmCxp11PNfe5Ik3LbUcb5G/hwItRvYDNBgQfKrQ3zmMJskWRPYLGUQvVKCu1cs
BVSUOZyw+UkwmwdGGn+KcJaFIu1fMZYj6t9SEudOBCPlmfVsXnVy2aEtunalc/U5
9sMPSrq+dICwtnGrI0MnLzBHqOqa5GAvHmoHcX6w04aGR/j9jyEFVU/25YiNxN45
QUGDpMNHiWS6NKDm8FPaNQS/ZO+SIXsxtKE0ty7ULAUJpQmCETlzipu13WQ/CSsy
WGIKXFKG4NjPeGRtYqCeshSYF7qnunLiVyFWknbkUA+QlbElCr5QJ0jNieKQdO1S
+7Zac9svHb3o7kmIIzwcaRGZDVgXRmxFeViBIxMAo/5QEdyfbZjVAVV1FRhA5k+2
PWEUf/e5qMQ0AtJFXwo1SLlOXb/1SO5zVfryGn995OiXNQWfn2wcsC3fbnUugIWf
+wi4ck7JQQAC63PydQCn1WcHvwzuXBAPVF89Y6HGz7hIxWU/aFlGiCngo9ATVp+Z
sGOEOFhY7ykRVuGle5lRZIODyQZxwDm7yLNR5ilQOZUGVgZ5SBXyH2jBngbRmiue
VyB8DLXW44y60OVMuvFSdOGquh/JsByVD+4aqATeBsa2JK8iC5+Y14ssPcZRpUj3
sgKY6bhG1Qkkb/JpDXQra3Mw92DRKg1lxcQBZ2PhfKeEYCKL5q2wxT/mq1RNdB//
jQN0lMXmH7OyIAYlv05MHnM1bI0QuMSduQhkis6JWlKvJutNUsZ1pkvsinZQ7wV8
7ndBL2ChSGg5PtlFxrknNfkLguSEkL1I20TqggWvHfGSnchRint8Y+wc/rQrw1T6
hkkd/Y52dvphV+kY7WGx0djM8GVfVjAbu/tJn63ofVqgnfoY6oKGXUAkzAYh2jM/
NQChG313HqFBfNwt+VSrUSSrYV4R+00x7W1QGlet1hC60xIrnCdJRGc8P0iIFhDT
AXYsxbH5ruNoF4sdmTZC2iPorkSZ9c3seceMQ24Eak98lJuMmk3o6P+IoipksvUK
1+au5fTft68/CDHdOkKbKOKwUjyI9vm6g43bDDVdWOkscJtot3menGldBMFhYKOk
82r4EmaMldgaAN1glywsF7FlNFoTBqNfjq6L14Lw0mgz7vOVVYWyPVhkFMCHC5xO
Nx5TKzSELpqj5P1qDeAk6NDEekSbI3NXRRe3l0nfIbG1k45I/bv5xmzoS57kW9UO
IcRaO/rR3Wm3g5yryZ5IxNDK1NZB7DpW+Sgm2+zCYLFDwWvslYWf88s2Ps/XzN6c
wo5gDiRzvRTmPyc7mg62QB+BK+ChpeS3IVqc1KdWutDtNF7/5DzmgpBoskJhWmTr
RQauSUubJ1qolf7us6fKg8Q9f8Oa43JtLv/qqDYtzPDy1d3qxfQCl9fSIbTHRVJ6
HSDyZgC2tSnolcDkWtWQtTtkov7v+GnUJDureF+/BIDPNT1fnLPVCLLPsHZJpEp6
HB3P1BDb4RykNO0M6my5goPZuwdPlvrVtuerJRQWfg9IuvSfYmdjJIVabIKZGm4L
NvnSOFU4XbG4rhHQJ1p1Y5/dxgv9Mirrk/c0dw/1cmZmLWO9SV5mks8D8t7HHmas
tILCdTZ4aWUA28g4cTU39YfO7WCbvva3D3n2q9+6G/02xLzjtqazUXcQqRYFedt6
fibgAwXy+wn18OQ9Up+mmvghdT6Gcve5Cls50XQHRXIEUl6P4Wf1y/kWHu80EZhv
K/oNDhhURefU8ouRR7+XU+Mv0a1LwW/YxLFD6UQtz7b1VUmMNHKz/W6xtaFXoqJ4
DtOc4MHiqnyRNDgcJBbDEk+12QG1MVu47whYBHXdlfROLxtwYXQ743KMuyyYoTMQ
9KH6CYoLxQFBYsOcNLbtvhnZmI1jGSl3b12flcqbt/lrmM9MWysOs6Cqlv+vbW0i
wdDJt7m7rYTur1mNvT112zI18BmQ8g0hD6OaKhp/MV2p/rG3icfPujA9CFxhGu9I
FmGB+5nW0uXTB6yiBBdHtq2xhPwI0++KYf6u43SP1fI0g5L7S4OX5m3IzgdOrDof
ei1i755RgGN24ja2RD4Izycc8DozU0lAQWj5vT/suODNlqRwu4IOJAAaMUsJWVNR
qTcFKZRkGCqw+GcwhR7JCfcq5EYt6r+uPhIfGQ9IRet2g6kVCiWp9ZgoJipA/UBK
WyqSw6qffSEHclaxCKEzs2v8X7t2v5SgXF6HW+ysKe4K1HvV57fjIkJb1qcqeXxA
7poYZWAO7Z6SS6faUDs0UEh0AJKyeCs9/1DLhQGWoUCmoGdFBpS2vqQdpGDT2wCX
qzl7xcXsq9nAG3b0ZUTilUHLlNVo9MJKeN1Qtb2EHGfIIifjuGpCBqSPJFTKbmf2
55S5t7ORL1+IDT76gahcTx3zTLnj4eey0b7Wprg+OCEUvI1BuBV7hS0w34SvdIYe
fsI/s8WH57UJ3S+sqmnF/woxaZOK6ILOfhUoNXXy3zU0qNLh6SgxLL+Edvpx1byL
5aCehG0vVs6m0U95LFy3ZlfbMKGGwpl7pkyz2IwueVm+OFM+1GhWeK1EIXfVn42U
T2GeLVT9m+KIYf96BgRjLTz+GiaTBvN+1cRbX0je7iNZxyYmgUeB78z+O4qfMC69
BFk3GAvm9si0Qys8GSCQ1c/L2e5KbSihQG8vdlxgYuQOU6kik0Q+ZZt8LZzP2kLO
XYxu+qKJgg3+7yeyMqbfg17U95muT1YMMJOzxFNnWCvWXdTTZe+qQUp8BRWAQdQs
b/kxC7z8exVAZh9D0NntGImWUT1lBc2zDIDg1tUev1w+vzwsxTunHfy9nJ4sDe1P
LLTftPKu2S6iX3YnajPEAWTfQNDhu5qS2kL+kLf5NzMvWSI4+FgAMswaOi39kNfa
zSMKEqQUagikxv2ah2OUqiBtGgkz40jruz55KKvQ9hGBUM3zvmnyf2jex0FazIBT
z1Vlzbns1MmPT2IBfib2+fb5lSgm4PAymRjIgg16b3BrD+zx5gk0X+g2OPDBjwFx
QafHrnJz0Zzc5GjInxUC6rSGnHfIBFdeE+WjOZKwAloqWh0DadgfUV6baTJ41nli
RxgRHPCQ0JKrzLdEDuAKh8NEUqLIYgzAZVePplIQAFULj1wc+1TVoXqiAL5Xh2Zl
HVcIQudzaUwo6Ohzpz/nQfu6nLelhaIRuGLyhNcm1zykyZOgrZDA7YyAs2jQPLNS
D3JZnzP/xPibKsmKxpkBwzetM+DckYneZKgu7Fu2KKL7S9/14/P5IMxSPSV+feIq
cyGZV2NDDhTbN1AxK6wwFUQ+ns/P9J0Et/yaF6/qR4mYGLR6eywV4U2RFQJYs0Ty
t5yuTSre1bIsMhPDu4jyc7KkN5U/OkkBb8i2WAJAhTAoWNv5TJ33p8qqvXIicCCi
bvFZi9YzMExPi4J+ivNA714GhNKHK/PPWoRSZ4zu7fTBYu40JFai5KPeW2+jXbRs
6ZeyPvA/0TJEQeHMlfe5kLn3rLjosGtLwuoa6LqJx/g1w56C6AGbrxJqwPpIs1Bl
cFNfGezNhOa/q//kQNtJwtmE3wEX542hq5mhGMQfJecLUJ+nxz7vkU6aTZ3HuMDZ
3Jp86BpQ2r07A8D9ZJsTXhlCVMG/SME5p0EBkVJHa5b+Awja2/psdnHb9N8LjSkz
nPuPqAuMWsm/YdOFJANP8FGa7RA0XNrGgasl6t6v4z4IXyiBn5U3ZEtMrdchnbBF
KX/31koaSr06SUeR/WPuwKH9mrW5WWQPTY5Iigoquc5ywePfC5gcNuZro7x1BDXF
BpqvLKwDHsSttRFrctxXqWNXBKN2E7jgOc+tcHjhMfqgvcn7VE55oWr1cdHmHtvm
+Rw9aoNS3SXj/xJaUqp7X5FjAlL7itumtX4Bdqi3Fxy5l/bymjMojcBbIpjmrKcs
LYO8N4CjhzwF4lPPSAA7ujvjIlOnwHM1MWBqlcAg8vKkDBgu3zHGj1+KNsWjhGvX
JJ0r69iKPk6erKH9r/u6IIfXK1RZcOe/dqtvalP1VI17Fv+7stSQwJpdJIwQidL0
DIRdnHfHJoU3aeynexVgY4OQSmgQa9agJ6rR9NZ8eBSuQj4rcOUVZqR2pJ5kknaE
gRc7o5hlWZehSUpCpjgX7mQ1Nwxc1np6AuArOGCJ34gVp/3WDc7+3vutPO7p7g7K
rijheq7mZ0PNKfa9CnJEqdAAn/Ow5kMULneqLuKC4zTqpNglQCCfXxRJdg9sRpOI
NQuE2Kr5Jm9MlAKHgcK6QCJlDXxPe3sNn6HYLNa4aIa97I+KOYH6mBtxVt8u+eIT
62m5TU6wPKSfZzm8vwM37WMx5GgXrQnnILihX1bWTwLUV8B5LNihuDgdXIQFLSR6
QCGL3U6kmC/WOljAXslI9pethl8rU/jApUnmvijW7n1jImhz1RXoMGhmNN85F1wg
U/XyEol5Vo+MywUUeK5y3evZNJJPAZC3iPZ5KX0sjcfah1DF/nbPX8WiG9NhW6PU
PC2oIvjEKeOyjEbGLUzbc8zxyNJbK1N5b90lzNZ4sYqpRWlLZ83jryfphlTF1s8Y
EHCFCuMBe3vW7rzvmgykjh7atFmRIAA6dtTXc7A2dQmZL1KzWpCf1yK21xrJhAsK
17rkJYy3C8D7zy/JUIyUj6n3mRXi9lI99XXppxDztHaRjzxc+fdnkexxlDlCEirW
sTU9dPqccyhM1st2I+FrNCuvsi9JuKuVus6YLNGT19d/+gMhkoD8KaMklq0fKsBj
8MzElC9VRc1JdX2X+59wgZ3ZhGINQ7Go8VKb4WbV1cBR2dCHjSvyPLTRUkRWrgoW
bNeV+gbwRmeWLc+wJItTNJhBB7mduMlCA1LrQBAxZi9ev0WlPzdHv3+Kf7aQADei
/f4a00kc32hQ3q2Xbx3xWKTO9UvxIumUnZVC+qS4G6u20/3xo6ckxhpDvURlow2g
BNjkzRNXSEoEGqJ8BmiXnCH/PtotM7QuzReyLtGtSKcmLR5VARNANFQWke2PK7da
`pragma protect end_protected
