// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
pgQ0EjONmfAA/fAj/lS0MAfyWaFFehOlFIwFSL5/r+Qclbn17/WeMhiJoxQVlPyCLY0Q3rnr2MED
aPg+vxZ8ObqEcH/9fcmKVkbBFB7SSA/cSEQFnbD82o7EMmKnSiUwwEx2BYdMwdZHeG4DmKcZAAfY
94D3iDkIR+PG9y0sA7xxxZqNk98U6guTFhVDI9Esgeyl8l293g4aHsUyqKGwhTGTxrI/w0zgzn7x
1V6EovrSGIBwnnHDnlKFZPD2+n1hnvPafa8AGajIgUA+ePuX+XaQV8rZP0HdQbZxBmEKTOx/WYu9
HjOfVijSYzyFeQR3SBiiAIcjp/aDeHcDXfYK4A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 13744)
mn1HaTAxRNn+AmgTuvjJTHqBcV7GN5UjPMvSIk9gegLP1hkhnmhl7top4MBkpPWurARj74/zs9/4
uA9lkvTOu38UMxCDt8J1Xk6GTMqbdb4ygzixFvUXK5C2NAupJMzu4DtFkxqyNm/A/z0WqzN8mNkn
7oNucfI5+4PluQ27YdVkTfMv2XKfN42MgCIiSfOTr4F1aG1vmrpZYzmDOg536lxFPzS9eGJINLKc
Vorr5XuRz0k7BncvfjKf2Dt1hBrn5fMoH3mhWSDp23qQSKAt1FIu76HZFRhJplCgpGQvZo85sYLH
h8p5QZ+L2C5LiOfMZ8Aeu+FZzisLZezQeGOSfxGPAuiPKJ4j46YCrw0mKGPWda9Wr0n3kF0PkqUJ
mww8uwgUrRuiQlscETDFifdVCQbs3CfKDAfvfHeGFpMPbKyCj3D7qZStSDCmzLhq1nzhEZ3jgyer
tC0+lm3a+zBQQpPH/j81uyBg+Uj8rqb7iwILL17VG2TXWWzu9gucTO/Gs8e55k5mg2zBqu9aSmos
wKzHQc+LgWDeFV62gU3Gr6gGWiBbn/WBtZcp4MV9iGSmhC8MfDCcka1pkzG79vpwaM+PSfZ+vR1A
DUdTlbxmSc9uowQ4PRqt/ZjQS8/u8KaLyZNUcQBreV3PD3VjLBW0p55TsVelVpa8R7hpOgEWCvYs
EwxBawmyshepv2evfZ3Rpyk/3uDQFZe/ZgCLk6fG3VUfH10MZVo7nLySypw623CDfEETLpdEXLnP
/8pUIfgFhmJ5GOl8z+JSMajYL+XR7epoMIe2Pw3mrikrE/Glc0/yHLvu65zR3BRpNqCFQ3UOqD9p
Kzm3IoOK2eD1AUmdjdgwzRqfPS5tN9OudwVF6S5RlyKMzSEXQObqOkBFFWkUEhfM5u84m9WkI/Ls
vIhpQP69HZmhB6L4/4mPl5qtpWnYW+4k6siAfzjyCsMI40+gsq8mFzkPFn0d7rLp0dQR8Se/PB0q
JnVy3BDynb7kC9wWMYtkhcMraMYoYnQi6LTen+lnnA2cW+zRuABoAJ7A/ltiZGaqhp3243iy6kjm
tmnl+qnR1mJ3sgB0aatG7nxkY1eg0SBUjMf1aQ/Lb7tdk8B//4d14Um/ZBNl94HuDwALPGsKLcWh
BswC8fThUs//gOFR/ucffukEjOo/+k2Xaznkd/MqmmROepnEkj1uAgncW3c1nSeY5g7GrnRfnjOV
FxeMuNxus67gmT7PAS1JA3tM6GFdV+XQ/5hQOwusaHL+4DWkxwmiuIHFjMKLSnBgeO3jvhamVuFp
t4/fD+t8ZWm+5sZ8PWOHJBTByrqty0n9R7bizo6oSMevb38tNIHZBVsA2/hyGI1c+WJT/Wm/+j1F
iezhZojjgDmmDKfPuiGwqOYjeqhJhOYSurqPXoV2KH4NKLkwfBlbeIeSAILooUZWgWoIH6iyEwZE
1KGacLOv5OFsa750Oj4dN58O8VaNUIa4RtrrPD9+RUr8SoBwXattSdZkxozyrqowaute8GgdTdIA
5opygNsWSKt8s+SdT9PU5Y1CSlVzOLaus0TEQhYvvznp62nll9XhBX5xBJIE0XLB0koGicLm4rt2
Ovc9qRLG6QGsnkF5BAftAKizPeDyQigacFrWi4bAF3cNOG3WOaUa7r8CqaTgj82C/T17/6DEwZ0X
fj1snCUqKKxalm5fupeB/Vos7e6hl1OCxYt+/VBAudhqIZ5kv8gpDEDUlOw3rUb4vWc8luXd4+u6
A8o9YCmVsg5FJtrLMBdnEkH8D7fvCYPpSAUfWyaUumRgp2nRpdkSakuyQWOyr84N6VndgO/fMyWl
Hx9eeV9y32bKpvFDhgq2R0eN8/v0ZJ8Oinp+wEdrCBXFe6S86IWbI2eUa3RGmVGwfguhur0JmIlM
qsqCUNJBg0SVLM5iPcgQMsZGqfyPsA2tcMeNWBUoqjM5ID2Z2ILLy3LS1ECL0CCU00cszR6Ayg/T
w2ohsUUz7DXlblzHzcSfPE940KH0xx/kKoLwul9zGiRwuVsUbjBQxVFtEAW38NwEa5X2RmkLB0r/
mXBHyGKwvOfCZzRIcGD2TIxy9LLLCRp4JC1ur3AnEKyz8NrBe2tha2LonCWXnDSt2X/SI3s3oDt4
MGIfWQJoOWLzSu9Ok1iW0+3l6PUKaaRA/QNy2Gimysy6qlVLCbzGhAMGsWjVQakrgftPHUiamqmb
MJGWbksiaPISOzWR5pbXnsS0uJ/Hh4bntIaj5yxM3lWSSw05E4bTO8qkD+iTzre0eJLqa4RFjtqC
V8v8denZ9FAWpzQHsb+8HABNBsNSp1trnWOmkGxWix1foT3v82g/z5OTYTIwf4czeOWpZAwbOPQJ
9KKnV2vsrsWIt3blz8jcMapi8N2p9zK63AoEQ8jj7+sZWmqRuvQCGex+ag5lP3UnUo7h0iTd2eKc
SKdcV1QND1I+EYlvyInVnHiB6jL7gsfyq9m5y/1vn2kN+4zhDxshTkumnVbLsMW27xN1DwPDJcGd
cizuqj/E9M1WTOmDFez9ryplitYDIsePCW/h+Kuaxpz6OFSOojw6lJB1kaCbbmtbq6GaU3cRQFhp
fn2DogVSzFHG00q9WLBdR7djal/+PtcCsFoTL1P5yw8r+MSDhU51cOWBjum00cqVRXzFh77Kf8bw
j1tKaGf+Fq4uSt4EjCgzmMQ3TzBwukAR/B32GQlxmLoqT8j8cvQhiBFVU2CmNjvIaweytWCSVgVO
o1wFMWgkbfKqNg+/zgryoh+WMgz+Do4yuBbons4Ciyv3dr7Sy5sjnvjVCAT/YIPaUVkEo5BfNpZH
GqCRQ3QFxijnp568ARUuc0LtgDcmMc7li8fRDDVs/T3+c23TjV1Zs1emKnNgp0gysHRvAlB66tpL
+DMCpNQyctb8oGoHDf3yOunQcUNDYk7Oy7eUs1X0BuaziiUpE1/yjeKgLa5QqD65OJUjXlkNIY3p
vAcY7jxJu1etV3f1cqgwdRAmkA7BJMkG/DOBFQ2Eec+7vek3/fM5hPvKMEbYK+uy9nC4e+aovHq2
wtpU/YJTxtyTiYQDj5tqNmomH6zOpP7VfpswMGKxkYVuGZ4F/Cy3H528zLZZdPNsc40OoS+XA+oZ
ABiv/+MiiiHsBxumTl+CKmXx11O39om9ShNoXQHvNQYb1xRmtFYCTLKhb2tw85wlPaKVvNx2XcWM
vEWABs++qBnvHVodYkMTmAAVvn2DsnTE9ugZNg/uUlEMJXT+Fq+xtGc55QYtMm4SXV/I6k7K3vNB
fbATs3/mSvM6YxNtuvH6j3x+XxNzLh43Xso6SA3ia5/PgE8oqpbpgO/nZKPnXghfv7acXtFe1ypK
WgQfb9M268DRRRns2jkxCYXU7XfgVZr6Qb0nRnyKNKSzb6mEbT2KnJD7KwQcmqXBQpXbURf0+V85
pqZWq72BOBsyosyN+Jw17hsjWZSoAJRqrwz1cDKl6wq3kFj8LFO3e0X0dJjnApJKmK5OTsBhyc0z
rWaQn3UyRUoHTlasNl9uOivBX2R15/W/lNmM+6CWfbrs66+f4p23H0XNEgYX2HoUJhZSLAYCCRFR
K5AOegsP92u9RbHVsB4VESavVq1mlUkm/0sp0BdFl2UVs5nlK9n30HDDPpbXF/o48QtpCS8qp4L5
kbtPeB2ofGNC+MX97xzi/aEadnp624sgFRX/+8n1Bn3SdREhasA0b/lS0Q5MoF0x0MhLcFXK14bp
h+LNxE+aTRfr5dnbzQSM1lzhvY//DnmaqnFpBjEf3kIcg+VA61oDtbvfrjafDWbjRSkghWiYs+LX
6kedAXzsbwyW9qAmcEflGvsbc24JAnZn32G5rkC5cHfTUSVBzGO0mAIFYeOlA3Pu9j+HW6xdERiQ
XmSScYYAezSuzPHKs8AdPUa0/ldrh7pNk4MZsnnykzO4+b+CvIS7NRCJ+b21ukmIYJqWb8hrk6Uf
aW++icLB4YasLEmDOQNC4y7V5uZvii9v7p8PuGzyRR/xItjd9wvSnMna4zJNcJ4cs2zuecr6Nuqu
c57Co96mOt+OFoKMraT/ElupNHdAiBz530hcWTDr/O6E6MV3CjFvmAo7lF/fWw+aecWX0HMnZ+NG
DoyZDiPh6EHJ+lcy2njCU7lkyRNODDPW+MYW8mC0jKKzpFpsO7JoIMtA9MEQA2J4k3VIGWC4D8YZ
XJ3AQ34LV3ZPty61jF9GMOc1GVFL8I5mxaTGZ4n92Wv2AXn1extqk16azuoE+1WP1r75O5N4ZJqd
q09BpOH8vu4ImJqHBRIEli7SHDudMh80LwToRPsl14rcusS0+q6TzvAv6E0+2w0xB4blJOZSs8UV
EhbkXY/F0WuW5eSUwz3ccYKSTEA+yHVwpxfQEaC90umRXvaV2Qsa6spwH78PIxNT06XdifcorHeD
xImND80LqV7Qx9uixRTiAPXRbHlhjZBT4fX3RiRfPhSIufgS6OsoOlQHCAZ27gh17oARMwcRgV0k
6ZsIMYhlYybQHB5HKWgdImJCMrE3zehn9wgxzyPEAFCuim6nEO2vZFkhvp3DU/DYUnTq5hlv0P4V
5aG8u4H/eMT23B6dd0MouTkqR11nADb3TjREChzEAKT7Z53ic6l4F/K1RAizWk0yb3AyxihwXKqh
hW3RUoWj/6jomozcRs/0EMu6i74/3+zgYb4fAsuafSCt/C5tcB6+Wip+rYiWcOpguyrbUaZ6D8Wl
a+Eee0bfip9ZYCJycDqL5OPPIIzgb8bNwMKKBfrZKlqyuhFAEECLXVyCzrEkAAAy633T0czyCAGc
exWotial5ucoGohMd23Wm6rFdI62zpx+m17MGo6Im0h/ElZa+OBxrQrtduw3t+yvb2/eX8O/uS1w
xJv5oedK8dNlFZKo9bTc/7cIGz8RZRR4f01nI2WwBir6V+IyMbZdXRAEVTwJpM39SA0UEd0J3nhu
Y62TfFRS94owGVa/36pYR2447gAcQpKI6wRcXvjvEnae8lDY3EC+NES1O3R6VlDZR7BsC1z16yBk
9kjuu+xvHIQ74HbnT5KMHM4qS8Z0vz53Rnzp5cSN7dmyF37rXMsdc9zkQXRLEKB11ov+WQMyDb4B
M56cXFttPB0qNHSidkLHmODl4kfUD9J38PFPWcbQ5rkKt7Pw1Oma/CagHRrcGcin0ieATJFCoPXA
4Q+n9IapWSWQW+LwgAtQrxcVBQT30AsWxrr4/3CY1KgYhStXI0dE7lUTJi0heD84ytMmRqca4ZL7
bRmou/68437LqGKDZuW/QjgadeU9wz8IGRZME4QfQNOy55gxhWRZhzwjx0aHvSiPpSn0O7KXmdyB
151U1+vUQm4+1T0gxTqKrw3YP2wxA5ZdB7/P+tAwhZKxz7LkrqDZOO4PsdSGmLegX+5GjNis/Dfe
Jmf+Zp6FDo4iRzlE0DE8EjHXXTuaYy2IGh54s1isn0kz97PW5w4Cjd2+RjibmJJoceeZkQ5ZIRKF
KR6GhaTMSJNFZ127eBXDG0RNIYBXd6dWQxaECB3/5B+926DZW7tAwOzHyqqWfnGrDbBEJjWVF/OS
Gw/JaxE3MOyXhIZfGc3/p+vf/CclCnKhRrvFHC1rz0HRUbA2em/80L/LwWjPAr3W3FLYwloZVaRr
aU2OaEgGii5vRBbL7pPf6ze3gBuXhAAW1XnGQIF6kA2FBz8pDrHkYecFG4C00TwlKlT4FQ0+Un2p
7r8ONWhCrNe0SPHOL3JFvCjooldWJekLssAp0mBw/nA6sEYqP3tUA+zLw5CKJeK7+qSmPjQ4GUF6
aleLZr3tqe3lC+SVcQYhM61UyDW3BFQaJqboF4Wf9k6/gz17Y5dBH4E/wOOrz4hYT0UK1fxwqyK1
ECOUIz9aeJvMa18C8mp/OlJBsTxvygbdzH3oEybr7Gn2gf1Yc9PQvJWrrT5KLi19Bg59vb7l3vmT
smQW+rpuPM00Y0QLYJECK5e6c+Iz+Kmv0kOFGJKazsqWl3kAovlKI9H+DyOFo6NqgD4RjvSeJT7/
AD8+qao5zxxqR9UFv5AU8zTJkD0/slWNRWWkVGcx6z8yYaoYD+pl/r3RwOAMJjq2Df8m/MRg1bwL
cAdsZtDMVmONHJQgFd2Po1R12QlAMDZWcUFzQLM8FjbjapokYGUWy7DNZelinh5niGdHqRJ6yxx7
VEGZXvCVSNXovrzmmhkBcAmmXK4wBop5hpE6sK9nmvSszmrK+yLLPOXkykLo0CincfH8n/SMWJKV
noyg02h+It4DVAb8b3lmDt04e5FbjVEdC0lym75Y+iuFzRCfR0CwjtU9ty5rkXCsqUHkDiIgp010
3jYJcpvcBNR8VNfKXZKAyOCqTr21sYK1tHiwc3/5/ku1qYFJyQdnxbOGF2tw16FxguadficElCU1
kXksIo5/JjUcZcWKZx/2qAf+92zwtX3pTgeKh52BiQ8g6QSjv/GlkrJi96KAeZKFqIjdR70o3azo
uUp8BIAkUdCxJF30Szf5ZgYTRZKLYl/Unx9RccNs1lKfBckMlO3iSvnOpsDaQGHqtrgC+xCtIQMC
+dBt+SnamR6kV/BQscSuOIXddOt9U6Ew0LXebmhH/87onrPhkCrm34UbKuazaI8nDp2+u5Jm+Ks1
XYfhnKpSIe5esHAHYXpHnIwHw64cCWx2vvQcl/WgkQCn19kVkStZJ8ufMXlPOFSRFPTIwbFR13UT
Q7fXdH7GYK+6IAscTpGX1zc0X9tJgNc1PS5JRaBHYA6MHhRPBq4VExCdbuZHrwbiow2dLe+4G+P8
MiVtdv6Ahii9Q0h+0JR5FB42/2LCmEFv+jUcK9hdUgbfMNI3fhhhh0PDPfAyleqwdekhDii8G+Wn
vuhLdHcgwRFnsCxLi5tOkQFAxA0MGUfcc8hhG3btfqj7ohltRq6oSP1XNUY1qk+PAtu9Ofe03Ew2
7p+/f6yfypxGpDahSWgBGZ9sYb1eTmxldrJ6PjukuWVUAH55mzI4nuSvUg2noYrcXXSYLasktRea
BJ/mt58gEJUiklJKQrFria+ecx8kgUQYvv6vg8o3BOuUnDjBMXt9OYkfvluHoEqjvdOXL0SbxVkh
qzGW87Tk6ER7WrVKMJAQXtHaofMJRwk8DJ04ZbRtE6DLtS6G39dWlWGS4SaGNQsUDjg/tRdhK3Lz
g0fM+0FIGH+VktS9nv/yEu9GNE0dpsUzOSeDhID7AKTnc6VuAF7vA9KKXQBnd2jkCiEBuI+nZV96
AHNrBvWKFN19j9dlGOnxHYeurO8dMCXuGZReU49BJHGOJTsWmnShexipWiWyWc+ZGHLWI7lU6Ao2
twS8ymIiEu880gTPaagWUjSMtdoGAGJHSpmTDFoc5nUch0zreObFw/Cef9Vqlzx+06UJgzG2UQOG
NfJr1p0XS920aEeF0IXilUpMhWI8RfwG96z0uTTPDe7og3oywy8B48hnVZW4oVYfK7XpuF0lmrjm
Zt8cokZn/iQayF6Zy/yD2YEm4QQ6v13Rr3BBqnrTlUYUeZy0YizL0Q/9FpL98TyNPUUxCX8TkdBx
T5RXsVxRsVolb0COa9c576InkdBK16evUcel/B24MS3iOfWe33uOeW1bB+lCKJjZjFF3MDWkYxME
mwAQTeChe1/duSWUmZXB4M3+hIlOEMuftfMvsujVn04vACS2pEO418+QvN/E5HfdOzNaAjrRjC7E
YaQFyg3EZTrmMfitpQCUkJNMfxd8lJJjoyXRJcaReWQ5joCO2oE/oxcJlXaiB68rOFHgmOSmCRhp
HUywvdrZVDdFoTzEqUJZ40ITUr+btFeh1rLBeTUQJVHnGb6QNcEELFfLxf3U2vTHeo+DKU6+3j9q
KPjQhM5CB/bXS2oXkXN1wt0gsXFSyCfdUS0aXEs190liGq0ScELvi5KmklgMKINsNoHRm/JWJpA0
D7TvirwiUBfCebsh9jTcRt1Wm0/hjJcuRJrRHTfqdS02xZyKEjEDwrZzz757o3zXDeCZIFVNOvaL
gYaL+Bw6trmqShf500CygDlaKVpDbrm93P/SbB4lFKThFZEaKQjBMeJsv74bhoBKOoH0HEb/f9PF
7jRAMed7vngnwOCCbyeYISjz/nAghV3YPETQgU/alclvs/2vQfCtjqbxDuJommhs/kISACt8V5kY
sbed935NdgR5Crj2FV4lSCG5IeA4uJ16zfnluVr70LYyen1U1/tFYgO51O8JVkgEk5ex+Xb5CTVC
8yMJr7uop1uHa6E0GSCAAFSAQUT6hDoQBgcbns/MVxLEOTfamaK1lgOjvB/q7zyKuLWvQi0Qj0C4
asN7sfGHoakKwaFXIRPtB6YRGsSdrHGg5KcvHHQ6Bbj9+WjQ2rfQiAsul5iYbi3OYQfU2quHIhQ2
q/1FUEULluuvAlnSYvDsYMVGMW+B/ttTSolyNwQp+CsjCD+cmXkoEHvSBDmmbRTFbS5Hr2eCwSrw
pBvwscyugPO8btk3s6+3uFN0SfPaU70eESSOGvz5HxzK4R9ClzRiF1BzRDxDdW+zANNQyhevNlzm
QmBMo2aTd2K9/aoOHVoibvyuqTvA5mJCOwSJSE8t2VYA9WbX2VSe/y/lS4kBL1YcMmch7KyAsvzf
XK6hU8DmGjyv6FANPNUFubzo2DSxV/K0bspD+EXyw+J9vb0YyKN1zJvw+GmzQiZuCCbvTt2ep8Bm
D5LKO70UAvVF1MClssUE1bVrSId9ZJLQTioPQZlmw811bKQ45H0iJ0aeh7adUduwx5SGWsGg/05N
pc+hnl3IzJuT2W2ZGgY1QASBmqRb8GXnQhOIK9x6ZA92j2BTaZqdl24ZhQiFfDyIl9DWZKPtTkz6
FXG3ZO3IOG+uq1w1xRputjmX91+SIfAz0jWUoAyMqH89nqM2T/rOmNzKmz4T+QDTm2K16SYDM4uN
5+PbqEoV/C+I7XAbhDE1DBAdma/gW962XOHY8jBPkTqe3THYX5YY0OSh/qklHiCqsdYPWA5rPkkc
BMJHlApzmrYFmIgW4SyxoKI94GS7V+/6Qp1CWRHLcKEbT75lVEbJNKxE6t1ftPb2vS+oxcbz4Vr8
MWLeWI1E9r77/sS4cXZBWwJCnzAD2o2PK6/KrWYWHvPRUyjsnT7P33ZFk21TGKtMcJcWXlfp/WNe
nDDLcOvF8ohWR2wlOk5YMeJFztRqW4r8sW6azezMrzSUKkVTJLp+VH85iJrrm5dtx1j2njUbkhXi
PV+uHo/Nmg0rJqqvQVnCSaawPNtKOAhrsyGNvOuhbLeIhaCgnPuiDByiH+40lHhN/OeO0tV5rWww
3aR22LIFdmQKuXT/yOtFe0MX0NBjpEab1nIVHA9LwZE3FCsZpiBPIB6g8YVcskRYgUT+o5JjId1a
tFnByMezusNGaEly5tPSfHV8iRj5tIBQf+nLQ6kcJIu/VsS3xlQhBy4Pmx+gSrKAru1LI6/o63Js
8J29Yp3JYfp8rkdwRR61Hm9b2Trt66Y3007nJuogHoruBXEM5OUP6wuqniOx4P0WIGF+x18CcvLf
XRNB49JLGJkYDB3rv8rGV3EC5UEbgd4f/holjH9YLRY2AcEJ/f/jsyHBrH9QHSM1hLtBFbvxDRF3
Pl7x+gKzlBWxu0Rm0aVi4uQO4hfcy28yDM/ySxRzBgoo3sxUcREO4znL03fzIsmyiR8hOulszpIL
7WHCCAVgS7ym0MX6rWid2QVTToQGW1fM49JBLxN02t0cS4JZMN40NnbX8wCS1sPmY3gR3lZMF9uL
NsWv5ldNOBFcMI5lpVlzAwiT565YHy0fQ219l4/E4whouVsSjbCk3phvO6muRarhQLL914XfTRc/
oVjG3d6P99NdyMM9Vh6DWzdRrI9IcQmOxp35pulIJuSglm3IYlQful6d3ppDsBTZRr4BiDknEFbq
r1pgllGpWSViZldm1vM7hMcz2TRQm7XhG5j2hY2A/Bs4mVnXxyFD/gfslwzZ/Yb/sfhmJSNHsMbH
XDcIXbkVyZMs3ZWD1XlH5weeqnLoX5kt1hFSM++gSzhPohutKm1CefqWdE7fXBvXUpoyKMzkfB0h
E0lgzjZuh4l3n5MqCoWoBsVO961TBXk4LZKdUNX1YN989SwhQEn+xGDuiHLeQ6BNMudSfv8LaL6R
g7trYRWMTZCJ31nTr2++tqAcMkDX9qEoZJVr0P0Q7btDbhBcZhd9NhhmRLw15rVHMONA7l6Wswil
e7YV0UWI4TGXgR1e0K9WnBTYzuwDW/2MdR0auIBJv1vHY/al9LTUu8hal4vrI1MgECvDjeIiz3tL
7NM1Vx+Ynf1r4mV1hKWM5Qs3+BGHz1XX69P+3RR1hHxMQVxV59zf3TUjPbfoyHBHifMjCa3xWEC2
P9F3n2pxkqMoboxtR/Hm6WsxvK4rQUUGDCzedanHBl4UV+j7XlDiKLVHrzmb/MUDzVKteKmoeqz7
s0nMn0uLUjzF2+pFm3omlxg01Gg5G7d4ZP5wFNYYNW4/JAvl0/1Uy3y7iQ9fdSHVRHuP5t6Riepp
MCrHl1hM4UpcVIsHy7mutdearFvOgexdS2DuC+JYfZxrnJSUZWUOSrzF44xrlmM4dF8famxYFKJc
XJ8hB/EItwgLBfZZU5kRiWjBlLYf4nkD78ZJ9CSMmd7rGMGL34lYnfHwTFAAhwiFpZm83/uCtI4c
xcBg5WhyrokYsmMYx7yc4lRJjNwjjBhRNCsDYpZDf03eE5HqVxjXpsHoowyunRQok9BtdTjw60No
duhGAuu1WOMpsTfEN1LCf56qYETFODu58RVfvA59UN7ivFgklDOJrCeH03laluC+VBDm08XoJVN1
8ZEqUexrW23OVE8fTSOfYhXhO2PQK6O7sOZJspJ9NMWp/JKX6H2Wq5o/LX4TneVhepj95I3sGMgb
URferI0mFUE/QifAbLGuZd8ay/FyMBXgha8LctSts0A4otTKg3GF3w4ySJkISBUIoKtTOsVoEXp/
w/67RH9TMLQghcKbBoF1b4vLqw9LPIrb16Fs/6XpWldT+c1wkQrBNlvPxXqmQl2Bl3CIdRed2lX+
e31pybG4OpYWENm/rSpHmOAexS/PGnnit5c9NEXG1ZpVTI0oBUQnTboj3JQRp35M0gsaXUPCdAVn
ZY1ngry/BXKB3Z48V2BAxpVVxarzwBHho347n7aNz5FB2YH6kvVmyJKxdUBwoy3aQF4zoM6gbjpW
nuUn5C+LWazg7VnRf0L/ZzOM/etg6JhXy3k8W90Feivev6rZUb/pt7NmWMdcbGLnMrAQQEMBsZcS
tfi29fWia7RBloUz02GZPMCWgP0Ti9oe5RnYm4Iyw4Kt61t64ChQeN/UbbkFp3NL4eFgWO8Lb8gv
DWFGkP8G1fOBwdvzc51mcaM+XqTQvmbvuJZ+Upczv1hEETL80f3Ts24wibkeOSU0rQN8AC1a/DPj
we1PfJ1Xqy/oCAqocnD2lDDtc/89GfXNw0Y/W5mQdLO2R6OcanjqoJ6RYfkZbZRgSRyTN7HaTIU0
mELAd9feYx1g7dw+gKZXs+ckDlyGJIGuYmGVqsf+FPW39A7IsDSe5xoGwzWo8iD3+BudVFMMlTvj
0zPN+7S7pVx5TzGKMfpTKusIxCn9iRkd4CiQewhFLnqJfAjR3o04gwHAe9fHDNYfAjlv9juoSwct
/0joigdzJtaUWtb5daKf11SevrpkKBDMt1xKQl0PA49hjuO7rj90R88908pIrklHAnPlG0kfc+uh
Polbhd+O03415/0PwQBDZXpXRMfqFdTBMubYzdMvaYVSG4QAx96oTaVc4yl/9iC26faFiDb5pcj4
rkJjoiODgQzOsKSnL3QVDgq9pZBYbdhsImmUsBgkawsaZLMQIibZBQ6aYuBwuBQ30K0n6Ly6XrLR
l3387MMGtzmNR+FegFsCYNHmypDOSqCJ+Vg9wLkORNeP9/KdTUkAj/aLE51rbJflTRHWVUJ9auL4
Do2Yfc4vrUUINW/AupD/GF/eVrlJfgVYTYCv/T5nxfC8A6wuYWraTexa8NdXlDDks0fLpIyt0+Ds
cIPZWubhZlDKcGOcLukSjMKbTk/J7ABC0EKOJsvOt5tO+WqRHwuwlF1KBwLmbWTR+vfkCVFm7IRG
SWzzuvSSZ2bBzdKXcNm501fS0amTFUQHXDKT2h6z4RcDk7FohDBgJXGkE4SS43O6osp56/B3muAA
OASltFqo5p5bBrXHAxMuKGh7/1GPiunioFUVdSBTuwqR0OmKzb9d4BX5ZGc6UJTmIR1Ni2uenPEN
rB0aXNysNXBd5vR/eshnOdosmyOLooUGBr0giOh/c8NMsJzmI1lmxgNmhjaZw7W9lFMppEn+zegk
DS9z81h8W2X8yWZFZ7m5wSkR8Vb+F7QBFkS9rX38pAkwbWJ5Lw2UV3vXkmz31znTxcV+YMCRTKKo
VHhaDahXGQKsZ81FQkprhq8b36Q0KyDJcj1I9AG/RjsHcWYlFpBYz/xVOiw9tKzUGHl8ou4kGj4T
TMEbLhTGrknsO3UQETP028PLGT0dE13tn/tZFuvGB/tbVyV+bsb6AEWB68+RIeEK9pAG+7RcUrU8
fGs239xlsnWEUqJ9Bp9dp5eAWUJfS1LD2usvUBfsNVss41WSu/+1nKmtww7DQdMDABhh2VxpF2X1
Ha4WFFO4UQhb9Zo+gQHZ5jw/ZNM0E/D61lrRVCW+52S/QfpMX62GRfoRykOIzpuQ+ln9uVvvfKUD
naoSg6byd8Gl9lhEvrHvkkBfJqo58SL8/lMXc/pHiE8eOZWlzjUmkBexE1gd+IDff386iKX1yDuc
dwFDC5kxV1wGvrywPFB90zr8qK+w9LMqraRyISv8+cl9jralciVgggLAw7nzD97y5aeCAI6hx/Kc
s/UeaoTiSeh0dQaq+UF5fcWgRHpLfHRL4L3FYMszbZIIr51VtuO59NgOnRxTpKswjfxskz1ky+yU
eZG/4OX/I2Y5m4kQGCa86RlqSCkFjqFZwsJFgCd464Ut2Rp3+Ecte9cMRbjiBjOFpcIExOvrTRSc
lNj7UddChaupsaar9rYiM19eruylHTtuxh86TL46au4jbHymrQCghzQpe80fBhbI3CgbnnLcnOHS
HoAy9e+eJ/qzxbDQdjZuTW6w1Xo5q7WwKHUqaVSgCGutwP8mPodvN2/r4mITP2Sg/ZRfqaLeb/Zn
yhRQVdjKXVIy0wH/2HkZDuRzkKWwJIefJ2uss58qh4TFlT7GQ+VS0RW5kchzh1Oo959NHQih96JF
eU+Ap/aGJaJEjVxAwfe6m+f8EzOWLpJEUNZsd3OAWZWocDVJVMOuGZmQGH8GNC7F1g28OiQI1tnE
fsJR0zEFSI/KbrAGM6NELKOxlFbxxJpy35VaMDOJ4pmDILfw+WgpkPkwqsrw0k4yHpxJGeLKUO8t
j+szFOwSxi4Q7qCGTihIpMLoQd49SK1u/147nSF0Bs/hzTxuOPOhf1qIAZIm+on6/NC5gW12Z+pU
LFIePT69e+7JHLTshzmq2qCSl25c4NAqSn+esRG9jyWXmBlUKeuGVTbsfXoE0UBAzF7Fqr9hN+Aa
BmuAtGLOQcwxYZiTQQEDz2bKaGuYGfh5ilfa8qK9ufTFQBAE8elyt6iqt2DNAz25GyzZj4U878Ku
Jjj3m7RYtuO+zy9JQjgbgIwAVj0thpyFZD6ZyPATavIEJ4SMXISIM4A9v68DpZDP8uzCCidtZ1v/
JRK81kk2r+jAh9NxmOjtBOvMe2BfawhdVwffLBhLg9WhgbEmXQsBcmPfHS5b44bpbzsfAxZoAvfr
0+AVGbweyOKvWpiAau7Kl4MDOxvoLbDcHIMGyg+3yl0lIQNyxTjyPxJmViinok7oNLFU/qgZS1on
ZzJGZc1oqVcXA3Dnqd9smA/7ie+uIPVaOSOnwbicXM/u5YUS3EcVapymBDt+iqshJFbBUYIKNB4s
LtMk9K6pvgZcYuvJtBzhFpWabZBWDX9dqBszoByi/KYr8l5RUZ9pnsyru8LU7o0DumMHVYHUT2j6
6DANndi9EeW5azEoDtbdv+8LgwCIr2pLHLV3PlpDu2egm+Wup0PTyWrLm9S0ubvwSv0SytwqOMOE
m7A2JTqLZ7CWTe4gPU01v/E9yy5KDjztoBg/Lg7rnktFZzQioBAL7avOipbXkJQ5zBRLMyB15Vo1
eaU7gDANAeBZQ5+6QDG1jb9vFS0eqxjTu8VNVCBdWVwf48qRmArAJQh+JNie1ri3ICQ2D7Z2pqnH
ucG4mygy0ICjVP0gU3TYO0zSr5AoWom7UB8zSl47y43caBpS4qGtYy8AxhBHo2Z1D9yswZAs7PEu
316dxnz8sPAsmWQF73P/1KxPWjKYDpsNCrY1BspIVJm5xSD+HySzNE2roQzY3VcXbD3I3UmXMw/b
cjUp3ZaEKMkwp50cGbKSSDHy+LOSKbLEbJXD/Yk6vb4O5v1IM0IUp8S71uA1MMUzQNFkK+eu2bRE
GO9Ims3BEiHfg6WWxplQJhVbG7pr7CBs0G4Sdqft1RNjhU9EexuZylLDVrL/ZhtnSTpL9GTkYe8Q
hxRS1BLf0bsAJYgi+AIyZBQGrbkMJc5ILypzqcYU5bM71DWRRb/aRJ3IOdchwBIbO3pKQKV7CjQR
vLvowa9+LdMaVokq1getS9QQ3WpAIIvmhh669HoM+sGqKuetDu11+cBr1ukWfSd0cWNf09Mi3AUZ
XKx4S1C5187mVvWYWpq461AYLmU346zaZA/egXbx1ahshlRKr3YitR158wy9cZ5dNe0EKbaVKxNd
M3+8jwb5aTOySWJtMT7mI7IxxAw7Pd2JGAVrqMQgEOOODgeRp5J042okqhM687/yRMjqRvetAI3c
Rrc55zsi88zW7wGLv70I2JZ/KpDnYrnGjGjZAGeBG2JN25wP8t9cGBAVGXt4HWOaMSMXUdkgzw2Z
DSnV3CMxhNKhg6i3ZAprFdsjQ6+V5f+t37S8A02TFFIv0RcF3h48aVajXEpg+TS5hNEOC5L7ySj8
KeAPlWInrHa4kWkdyYdL73fksZvP0gXpv92+ICl0MtiFqn+cmISXirU1w875AcwwQ7FiKeeF5/5s
emhfL+EM3+4rOkwm8VzOfzV8sP4uYtSP7SmvV9Nwfsn8kvgO9bhM6R//nKBV0eseGNgEfrVE90Vi
Aa7vsGUEqI5Gb/HbG/6wjcolWbAdm3TQYlJBIUGNBqwXlNYqbN2ilcxU4YodSK1El2qRNvVgy8ne
X/mP8piNqfGN4/LDh0RiqkvS7wcRJYD0MuiN0g6PrmFKjTTuh9f1BVrIklwbF8+vM+pfR76uq8JH
F9n/p5TvAEafUso+wsC0Ugax0GC2mWflif8C2kzEhxMYTsGkt1U+FqDJQ84hYuz1ipWrOQHm7PWr
EcGr4bViFWvb9fT4UzNTIyIDhFX5AC1D3/r8l9fr1QwL4fMOBsjrj1pgS8h23WSOJaHibzVYrF2E
oVHVEss+8ntQIrK4J1JD2MK35DGGneU0ERLB+J0EawfCRA3CNfTbzHB3fQRg+zDlIcd1AG+n79XU
HCQk8QEnwB2HH1ayiWyEsu/CByIe5OuffDELmTGpXqjI4LBt/Z/ACmeXyM46jppGgDR30A1bbJST
mKTdqH3LCQq4IZzQ0KP9hJIZcVC7xlOnaHq6p4Uq/rgoQ7fKcNypWv6+bqugjglQc0MG49ih6Wz3
RCybLuX8jYpK3t6IYVCRcuPMNiZn6PllgrnskHsEKNH4V0G7p3Mt5otd/8Jq7tPGhynBc9V+AyaG
eS0BXGVLdix+kBoD4Rr5lLphh0MlG7crpqJjBa44+2qg0d3h2jo5g9dIDnOyBp6qDeU5cNXGtZ2c
ZcR5IUhSotKL/zsqSRPY/CQZ5N1HoJ736ULJGAKBEtoABuz9CSc+fn7rZOfmCltkKrg2FTqLgEtd
YPtGo+RwWIrdkFSN444ArGb4Ax42lDYvpFc2an5XlaseD02RgSG9OyE7gdXPZYY1uRmotOt3vuvs
XW3RE+G6SauRPjBHrp7r8CvUs6C/igxggvploYciQMDzqF3ll4Jcb35pYTxfgfYAATROZzH4kyT+
vke4tlZxX40jE4Yjw29q9ucoq2DQYMM7nLfangTqamRtqMXm4ushquqaaJWHGkfTUHix0Kr5/QD1
mMohbJ9Jz/eXlCEZC6MT2g9Fs7iXscaG/gvYrNd4kC1NUHR2bBPZ0uDTEi4MRvc3w0NY+enowSFO
N3n4Yfnf69iL+tW+2eyAB3VMUzlLtuQ9SPB1xs3OvK6bpdCIo5pIy+RrTbFykfE5fHd8+jJd9Ax/
r8B7WtpNsWTILwhC3hxUNvlGmRjccuZypFvdcb4HyX1ptkuACSVilvHm6QmEA92DRtajQtpl9MxH
qqkJ1xdK8g/rFJ3TPzHBGZLHufMcW/UY7czMS6UzHYTltwyeoCcSmnRoL79iqeLidvMjl4MA0YP4
q8DMXVVyERAAZRR9HYZtywHc/UmJJ9JUqBkPn2ZMQWv8eWk9fpi37IZ4ZHfH6jL3aS2u7vq0oq//
BhJfSQoCO6tNLuHvjI12DASNmsUCtDTqyPpseOhWCwVibPvliXtpoMJFfQCO4MIBLMXuLJdFWBnn
z4PTLfqQPy0Tfe9BXQb+FO1elC/fgJmDSFITGyF3vZVxA3CnSDEAfT26M1QC9HRqq1UQ/oqcTvcu
C3NnpRnxHpP/j29pbkNdiXBZJNmxX01lXO9laivjax6LkXNJKy2KvSaHdCa5KGRPwY/o2VGHeCtN
VbS3ncfwh81w+byi6cvcZhBiOGbAIFxRA3NStc07jZ28GLL8oGSI4ZNrkZ76s//GU5BwW5Veo4Gk
hiMiycBlhRUoU7ptYOcKDB2HQWc5z+pcy449WDtjEbJUzGB8EswW6A7MgI9teyuP/p5V1SzC+dx+
nQPA6Kb65U90WOR/IZ1wEm8++mtEXthFlqoWIZS2eL+KmCHQMLiH+aWL8P9FwBfXuGDjOt1VvomW
IQsWJiXvYJ+Fov1H4NOkFtgEyYBwEY0XnQMOkmoGGsbk3AfS6NMbAqWF0WiSjllUw3hcwDUxBhxN
bAyb1P0HUpNbcj5svmvf9TrjZ5hg5w0NBhIynPTb2qWsMCfOoeSKrnw46fmWf2p8Zwnf+Sb750HW
Lekx/OuFsjGErwwSc8UyYdIs7U9jfK1Jl7lw/yBtt7EYVv90ggNXKn1nXnR/wzWyfpUBX+jeIRUM
mA/REci+XE4r+7+hFoguHmc4dmat/3LTDbG0j3T2LwwuEIxPV9YauAFtUTIh1GtmCEwoSdh50F14
uEarE/rHXLda1d8YpzfUfS6GtAvszE+2NbdPUJpSkGzbqAtRYkRsyKgXw01BPTCWDjWz4LRc+QUs
OpWVkzADdeb+yocgnUzgLqBttOyYul18sKzam9fLST2BgIneU9X42GWfyzyF3rz5uxghf6hkuWl5
5tRB15quDTo55oTKvOz1F8yxcYwhDtB8U54QJYxLifFAFy1H8dVsJI8yk3OjaYeyqC2zxw8yHzaJ
BPDqqpB6InqhiHPIoApTCXcArZ/sfXYqGE+zQEUYXX0JoT3eW+gwm14cj+RpwSAjLY68sUl4m7pm
Acrs6bKEhMAvDe9DF4QbUoq/0h8rhpKqx+wWXXdkAkpc/TSgXbBP1oTg0FBan64OOWdUtdYmCAqE
RiNz8BYn0KjP2wbHbFZY+SHv4Q/ntYSBpQA9rGRpi5LB+QptIV2B/Q4g2v0WC0fXU7GKq4/72udB
tFJwCHY+0mFteoWtNh8NiGr9pf3L1rN2lE3sz26Ly6uG6lAd0D0iERTranYY1nDeCERDG9b/fw8o
XERpL1+Nv1Jbx/8NGKW6QiJhnYhUsD5tyKI4Rs7VaM6cqcx/n4jlqcNg0mW8hx3wQrl7r5JgkVeU
Eaxs9fPkcb0XpYZi57zmA4e6twQf+dWiuc9NEwuYc3QsV96RyZeUgEv7lQCvO4arQrsL+iQBXVxs
I884JGIQSxbURDXjuvbTPupP4/788If1SWE+DlbuPVp9cc5PNORyBbcVTM4oEioaD/0rGbEFGqp/
4lYjbkWQReiRAOmn0SNHuEXPT8QejbQc4kTEfVt6ZUwnKvdgQEsF1tCCWgx0WzCWFSVdbc56VC93
BaTdhOm6reGUffp6Yxossc7y3w7+VQ86pRR6K8wReZhci/Bt7oAbYiFzcF2lFPMubSQF0k2xY2E+
gDQdVzL7wObxHv91gFZRx2mmUbCybRORLQVKUXze7s8hrOxAK+Qj33uLWdUEDNNLfq+zETewtEDJ
KXgtrQpglAchi42891ApDbS+TCzNq2oFXXP0Z8jVwDWXt/++8Pi9uL76A56FviBbMbR9pg4kDscK
FDwcqRgtKA==
`pragma protect end_protected
