// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
I4vkCAAuBOpik9GdTllDgLKOldvsHZysWAWr7NuOFwN4widu6weWuo9Xm/SqOPBhrUjtWqCr2mcY
pPNa6hxcPFMBLxZgxoy2+jG/L7GI2h/Vb/ipeUcd0ARcizNuuICZssaqZe0t8C3fDR2pUkZopTLR
C9ucAYwAl9Qd3oL2uy8WDlmEs39FJkaGma/MFS2piMP9CQKMLD8XhwwNt92VsK4GuxNCNKnLDl8J
/SYHYVo46pFTEw73P39NFFgXAoTQPiDBbYu1b/4nXPXwbN+KqUP0DGLCiLaj9hrrQKvjE31Oakpc
HDDOiniM45pSWNK8ZsAIXIurXel7/0KmffLyhA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 107648)
FW0wxf78zWs2X3pvKeb67OY524mAv0G1HmLZLGPKxfGrnyp4th96GcfhhNNQQoB5Lqc0K7VMC/D9
Q++WYE+LkOdCgw+DzI4to/Bml09S5G1/86zwGAZPIzXrIW4pOSkyVP+Tc1HSOQEJ1wq5YUX0H6qt
bWSCfLJ8bR1C6X4s/BRrPVNuXLKa+NtDgwdLKW/bTebG8VkQQMH3mNX/spNzbMY9Ddo1Y8Wm7t7S
x9dnNt2DfIM3E9B4CqOvYJrp6Ujd7fryN/76zcEhQpSFbtjlwxmFeEC/CD0mOUGc54qjQl0IpWtE
kqmyr6zLCrpdnln/JzEfrhZiC6WZFGkSawUCHF6F+HWHOuMUY1Jw2NqIARiCIYJs6ulwBjR93qYc
nRfh5Rnc6MOm7hNOSeoNddkMHkDRz3TRCkQIv+YdD8ycGC0AyL4tyFBkIN42q+wpLiAiADJMkfoz
KGFZUv29x/TbKXuVEwKS75MZeWNhhTO84RhCQx3w7WpQ5u10MAgGKOFL/IdZy8+3wq1EepmDNAbs
sj5w5LavzKsscp6OWgTJcHBH3xMAZbXqlApcQoqUeAP09MVMDshG2ZwQSGB5oh462WyY03K4+4rf
LxOBZl3CiUI0g6jmp9/rSo56AORPolwEuGfLaazBCAyE4DqupScwoyYNbVkKt1y4Y7Z6qg3Ny9Dd
+DFHHCtnvoWIBZ/pTPqEJU7dp4n5trQFDHe+6Y4sP4sdF+fkz3hsctrfoqckah9czOewzti1pxfR
R6v/fJ+/2jN90749oOXrWawBAkRlnVblmsm4nO23SVo9UvNc1dZ4WJyvfI+8pRG+M5DmAQsgxnO8
mwsPutHjn6MhH7YkRSoo4i0/mHQKuAO6g4sy9ecHy+ybTUz24uqL/Rm/6QVsXDuPl6YCYJ8dIFP7
fdPhS/SVjmuQBbof3+vxA/XQZW2tihMyBUmIm2t3tKenAMb2PYrSSJmGxtFksUHL/JIERyLoFikC
HWXA3aeB1+HZHkgG+/o4B1czocvObfURctl3odoOX6jjnpaVRHdie+2P8MEPRZ+uPVch1aI7JsQh
xhHk63zqW4h26CY00Xky7b3GqYQHa8ZQ3K//CHQCT2VIUXSvN6Hl+dR52iSSuKu4QO0awMypVXmf
vLU9rzhFHZENb3Z43EAg4UduIoFhmPnROsOgL9XkbNiGa/+/sewGgvmnGyNsu74PLYBIfavqkren
St4N6peP4NmkRZvhMyPHDka4WJyWTdQp4tpt64twljC1XTDV6sJYcsjWg1fz2A10H4LCDjJMEeRW
6uKG8ymA/35kIGmmU8hmVLN9lJ2IziDVEt2bnHVnKOtfe+2fWlpU9KWn03UZ1IJBvdHkl7N8n5Oi
rLNoB/JzvUpxn4nBejlTFX8GmVZHLkxFCGd8rSumuKShcKkasW1ruXnesZCdSaajnQtmDkJ7NLJy
Vle2s2qMOVaAtkiDAHcZyCglUS2i+IYKgdgmYDPMYWfyiRwFp/654YUM4ZgCdTudZA/fHkJIHo0R
06eHSuZtXmChWRUbrVLwzIGAK9/Qhn5tsMIRYfv3j8cFqdMSr4CjFWtk5cRBhty1UWBPWHKxpJIt
uW0DJLH8zsGqLdmOmBy89EmvHQTrIt5bdbJBCWacKUfVwjHlA9KYWuov+kojOXGcYj8gqILalVd6
FoUoyby7m1bcd4TmLsumtM6n2Cm8VE4KSEYxEKcvorMVF/S2ygUyJczq1kErcdPoDRWBMmq0sAEH
JAuTmiTH1moHLGPRF7119Ou0kavVQ5nhGQ+8Q/QqJ2qregkDkdS6KpQ/ydUa5SiAPzVLvU8lP4dX
Drf3kUv0BPoS+JsZeY0XR/qmzXS0e1G8soRx0v22+UEWLIe4D+NyAOqHiwzMPgwy8N9yFZI8fFjR
TYG254ZNoUrZtA8FxQGnCy2tPE7Ep9BEeOIO+ZLs1WXPX3c74ZIJ6dVZTLcBndmAukyI4ODlXy40
6MQ+jF6OT7b4QhjfnfJ9hvs2QJrsabPXjnBnI+A5bFNWLpKhNnzP/UuOxwHJzQym3gc3fP7Fwvzq
5TvD1b9TkSStan93JqC1y344XgS3Ro5BOrvFT5N95iDUJtW9oOMPY4P/eECW7717JLmxHQ/Hjfan
QGMid2j9ffIaBNC+6YZfITs2Yri9hYztKXqm1nHFsQVSCO3u0veJWT8ZKi4sFHNVS1YKL4KHeRjR
nuX+0omBjQzMXWPEWwUrt6M1ZJ1sKFRsg2TwFtuMWxcp3ABPAggrFfHBDijFGR+LFkoS73EQIpYu
uA7KmYtySWwKXdteZFdPKCKkHbjiHq6/YzM+UUIZTSeCBqtMgEPds9fnNwwiYihaPleL6tsxBK22
t54NMLpOpSJ4GdSSpft5v9hRAy7Vva6Wit4zQAJOqbAPu18gtxCsqQuKcjHFGIb6Svkn5+Cl8f0b
oxgpb1RUJMo/nGpRHqABe83VsyEgm5Dyq5yPahJEnAj/XTjCml86VovNWBXF575F/CVZnlOK6tDt
HMytVHq9yq7Sz8EdH8tpMa30cY0x6A5YKUfn3wzksBDwHmB4QWumOtc5k6A2X9QqP3pYNLWIM6Qh
FoUfuG9ChYI2zyqHU3w1rA8qCP1gkLfYBXcNQsKUfANAnllCQudaaHiS6ne4iIR7D30Z3ox355A7
g1uPRiLOwdqYFnLphhdioRh22v2ueIVrLh+3JqAsY2pqyvGD4aEEwr7bALwg/DGAe79oyrXaA/QI
dQSF7V5VNSQE+fdn9s/1w4WZ3ewao7K/u9kkpW6S8ffimi/RJ8SrdztDIrl4gJWD4T7DQW6/B89M
hEvvUD2wjmJkiPY1iZ5C+zZtU1VuQOXerekuHtxr3VQiIDeXeuF4qXSdC42UAF+jCiC1Np3iok64
5yBYoIVLtCFhydTSldmqjzO/DIwx1E6ks57Ogqf6nFZQIpVSTaI9+H0VtwgsDbxKKIGhEmVfk7cG
sLH0TtYH3xTqpuJkuXoKItzBu1zpcCLaFRF27XuVbINk38Bc4mYlQMp1fhHY+aowyx53S5KjWSQN
KnwDMzr5J/joQon+si4Ou4nlPEl7c1at/Kxcy+qskWHh3jA/s0YDBzQckhZflpDNDjPeQ03A3xqu
57kz477dJ3ETWxQaR0w0b/KaLFSMrZASQ9HCzMVPqO+oGDON2JEUgYzcw9R7PStliP2/Mx437ztZ
f6m1Dxt3E0quWdRvw+1OtqNKPMbIGBXwgu+gsMoiR1AINYGw+hwS7DakzH3UcpI2z/Qp6+DVALwi
lhRMYxYXoC7tz81mvtGPp4nxtPfPNzaoQcWfxYgWoyammjY6BZyA/ng648IuhwUz7yRBHbSkNThX
xcQ2J2Ym2K9MxLiRjsjiLak8/L2Pj5stQafBDk015WiQCsyGML8M9Ntt4rDJ1URfuJ244vRfaC+l
RHFf5NdfRTyw00DUT6Ar0iVun09UkGGqCht/i/+mb4gAczHDrwnwcowc3jAzhfgAghfSd89ZeJbx
KCRMnQ3P9A+dEXZGwftr+LYCr4AOXaJBeh7pZUoEv9VGKiIZtEbraW4a6nsKU9GIlJtjiv3wbfw+
rUb8s0j6ft+nbGY9PPMaIFurRlSVf30wse8sP1Ozjo7G7qqJtA7Zhcuiuaywq6CGc4POzTRwp71N
m2Yi8lTz/WCBti0yYc5ENAwTAWH92NAUZj4VDbZtYQ4wKZA0UN2171KyRABK6x68T/4s4Gg0yCbJ
0GbAfgVBLszNg+2y+B/jI8gpUOGf5qQ5d9N1QULCVt7kMiPaSPAWh/Zug6w824ocny7IR4weHQCW
Wt5irB+TCVHkAVyAZGzov6ryroIu/Qaht2GcqwXihEB2OMO5wZM8Xxlc1ur/ahlFjqCsVzw0Oiwv
i7z5feGvn4h0zQ8SVBAQRaKNcXUZWowEvdnFzGl7SYGQg3gzAtzjTcQpvgL7EOlhgOJSBPY1uRst
XO9z8HdrlBjyE82oypJ7AM/vj89lSQX9tZ/60UkOKBzweU9ZgHLc8Iw/TgHYElY/eILCP5Bu2QNd
UnZQ+CyY0zVuMNkko5uWNYN2EXgTyTkvnTm9KfgONA3WF8Fidd5CFwFOviYVKiQeCCB5XfwyHSty
mMJtmIXEavDn8TRxCYaq6yqDruZlbssXnZdEuLRGl7A5/sferBBjM2AQufx4HVi3aRvas+UyfZhs
pXvUumM0L9K1nk7gKm28o0QdjXmzvn1g1mjVeMCGMGuhz5xIAIkI0Icl7XbRfn3uLI3+vp+wOhN+
FzSY0PmP8oCOn4Khyp5uBffPvJFE1l5biw3FL1Q9ZeNVdw0AahWs3A9MTr/gviig/24nAihGYFLL
8hdi+gzKgfh3Y01jqRK6sXS/0hcS/zrbw81zrzmduTU7dwm7oB86R3+BqyFcwD0yULrM0yPCqp2S
G+KU0E8YR21iwYpeEfg7fp8UwdJ5difcrgABnQTNrX6GC6VZnHjLb2/+ic0htNLEF/1g+JVF5cXs
FzTTvVBkSn6Oo5XzKT/ZX0fMcw5gZSwfMw4A6JkkymV64jszw3qLtomLdnzoCyRid31I+6pJDcpr
zUaxSh+H7REu0tNDwbZ1pNwnrIlIaXU17LfnEnvHAtZWKJgnCuqQb6igbF0r+3JJFaB9sqxhwx8i
E+WnmcbblahAeU+o7Q/1Dv3ipKC9qu8AFo+X61JvngKyn6hJW34+Q1dp7NsdPLqbvGurJ2srhTqs
FqZ2qWdrvqDMjn2Kn4xpABkwVrZLBRYWxLfrZ/ZeIxxSQpzXJuH71TgkrV3n5BfXJwMPkhajBG0O
zafj1ltSdxJKIDj/Q5utpRJUOZpJGqZRlxo/7y0MMlx1guBBELrz/IV4tWYxA71rVmKif2joYj4F
n82jFYDwvzQTw4NmYeyM304zErsetlb7UOMhSIZo2cCqyeOssNUMi8LeC4lBrC4BKvwl4UmLR6Ng
GY/seAawwY/c8nnjGNfHE46Kolnslj385kWQR9//RtuGlU7G3ZTRoPEvsmdKwtp2aDbr1Cz7A09R
xzRgQbdxopIYZ+P1HR9OaY1T27Xb834pB1bfxODcW6tnpDMe1s+14hKtW49W8bOprtYIJ+LjiteE
f1oRiYlBWzAEZy8auF7IZ+eoDhJBZCXU9Kz+w9WG5PjczVHNgTMycdB0aif1IoM5K12/VV9ujPIt
UpcpVGc+DppTJDREr618bUqMb8aia732gd3E6KrxuJl4HjSYxh4olpWQPNuad/Rzu2JNF2oRD9yj
qBSFW7eCXBrLvjtEYSrsg8tsOjUVgr6c5KM8MevyUS7IOcdgI5LrVbtd6AwcRfPrtohuzsoKFGSO
TzY2MHARxpbxVvVFugnbbK6Go1KQzJ3E9r3bYfNquCNwM/gzTPKiAWa/shFgiKzRwDM9GjkjvEKA
u51vr4FkLXuzthjld5XRgAv/tuV/mNbtvgBSU+/oOz6xyX0HDNiAMRDSfz6cXOZlXhOCcqZow8eD
5DfZ++k9SogV0Z4WnVmQ7Jm9u7etyLQvb9KPPOZwhMP5iEco4h2Sm9d6tEG84jagLGEiQlP6vaOv
f6Erebvry3CqYo25UCfRHwcZSJoo/SjMR2y7OjVnS0ai1pWlEXiYBqEC9O5wG4m6dT50K+Mf0G9X
YOmjmDfe6btUw7VF/h2CbJPPmP2uqOpD2yC+4GmI3yg1IQX2AfllHbxojjL3AdV90RKMOMexQRhb
D6rtme+8ozv7og7lmat177rXsZZl0oZGr+JbqDHHZGhZLBnWOtM9oMReQLMkJWRwg7PTEMsIkfj7
5+P8vhUOh+ft3VC3vx49gaGh5+xZQTCL9k9GgjKh23sNnLuo9Lx5BjDnU9ie+Sbqa8cBCXsl9efZ
XXMmpRhB74MpY9g61i9mi9BbJLxAOwyV1QoBiyhqoQamjMELxcsxqdvgXKDMnlBJKS59x7+aGyj5
2tcOixFbM60afULkrBb332bxFCr+SE1QlLLCfBKR1CI23DQCz3/nflFYCpFh8uQPvHu+WbSaOTsj
163DJ4QaLqMZqz1s874vf8YIsT2H+9+Jt4einhSJFZnISVdrJSJ7bNTcVxD6/scs06HJHlxFSkJ/
Dt3UbGRYNaU6rzDtm/uzpJylrkjQW3ZrGGnuVbOmbx0znJr7YzMUtbJ+Qs+1JViGOVPEGMxapIQi
SqGgWrs+ULTCnDKO4wo98mHljXREJeeg/cJSd5IBshkTwuB1+8bMdkKONTZJAwAL9Ot3yF9Z7oUK
aLUaGWnhqSxE8r3wG4t4Fbg5EBMVL/b0h3D3zRcGgSL5MiejsuDcMk9azW2KpKb/N8vADLVKyhff
mxR7+UNUjMSh34dY7RrSp4cQWLZ07+gx9QeY8RfsXgFBeTKHrQ7KmtLL+68zKnQVNV8qHbjvhZET
9GXTubn7fZT9r4MJSBbuA8xNN1Xz8U16b8yHI4wN/8TNuica9kNDlXPFD0+YjZhUyyicg+TI4792
ehaKDzm3tg7d94zAg2EiWZhoepNXlQsEhlPh0A4TMshWcA6LvpFw6B9jg8dbn8TH1hwHR2cPXIAO
xj4nqbNo9mipjONjAfxp9eQUzppJwnQor35o+r9qPvFcCkWavSUB6UmVqPztC9R3HkFW461GKLAI
uNxb6jo9immDWYguKv0hFei2nMynGirzXd3VhR05HpvA7RmZBoI6hGFN41HvIaxmbq6pA5ZypWpk
C/1BHR+ibXpcFDNN2nBXrB+wzDnotljony/DXMedv2Mj8ASDWnD+nNUQiV9vvqN8f0IZCBhjRZJv
236MJ6HcyqzYLd5nazXb/QCbKX6hfdZqiaz2vO5RHxQ/OmGv6OtxRqP3rfyIi6KyNTUmg14GGvo9
upaS+9Ck4RdsZdHA2R0RqHEifnCipS21trAKaAT+MVLT8YOv/mvVB8kj80IOCCOsR2q/ioIQDTO9
2FUanQvK+l4P4YtlOEzu3LogU3oYvsaUd6c2idMitW1TDIj9ryaZfYRTpDxM9YcoYq1UEBsoeVzz
cfTrWG9yvFlkILeL682BScHefY0KGMOZjAF8UULoUhKMTNh5kkolXGHDV4+T4sRsxT+qwFfHbRE/
hZdh/LEIaKkg6hJLcbe5/lEVBVySBSFMWFMZm9yxV3H5/b2ktQKj/y1tqaBmWWxrmGASiS7u1J3H
IqCRXzZ8HP1Ly4Xh213F0BCW6xjIazwboFcnfgVI6/8O6OU0q80gzy/KkjxEIB2H2RkrfMmHH/4d
fiU/JRS95SZon9l2UKaStV+zxcHdkwMrs4bVjs09raYraJDIfTrdkpvnC/DBJ0Z1r5CMsUMG89By
WXLIJbSF0CZFJhdAgTcs3WFCWLwwBbA1oqrp/RfqA+B+aOb2G1g566WFnYFuCTqzkyHjEH1RHuwS
hyPTACFX06msel15ObNpfl5s5ZwgubHEsRnFplWYEdj4Ar7zkFdhZ8wOd7dp0oDDvwWKzbEidJIp
vxuc/phM3ySLP4EYhA4Aa2nADyHM/HWf3TdV+zC2SLV2U/msnsNF25ruv/1Soqv/ZBMvFzRdjFoW
zKzuXeiELctOSUw+VeEufxMXkzA9Zdqaazl03r+Yp7RvLjd6TGlQkFUV5L/MisxXCdZqnjxEz21H
09KUbgd3xaEIT9lcpPRGpHK4a4BHTI/SaZcoJixV9H9LKP8fuZ8oL0M+nAuIgPIB9rTxTvZJGeEm
ILNpnIzJVI03FVlwujYrNsH0mqWolPbBE1VNcWTXmzwGze1gjd6X7C0wlSwmZPOQj+WdX3d/TSb/
ovJ9o6D1uZBcke4i0SW/esBE2KrzJSxRn+mhhoft5YD2szqNlUb+nM6XY664OsJlVZZ5dCzeXcyR
wsGRdpd0+N2jgrjeH0iaHccLWfQuFS8AgRSYkBuBtUH9Kplw9tve08RVKt4iKL0tDHTTQea5WG5y
HgILEXwdhDebjhbSWoS9Wz8U9ENaOtbDbB+TQ4mG9YJ7YBF/aAXA2YsbWhWnl7epQbBlYvINZd3U
i7H6YJAsGmBw9dJfvIp3BkwjOSgSD93b+QeMZ60PbyVm+Y+XcBylj8V+YtzqOY3LjpRyBIMeRg45
B+3dCgYZkQGPOzLpHoFGaEoUXJKGznv9udZeAUqjioN72fjoZ/gG8Gb985frnKwTsCjO+nVsr7p/
SGslOBp1MwxgdEOUHh7UI1ZKv70LCD9PUEc1M5Ac9k87pVVRNItQSwatC/clC8O8Na4Xu9zJObnS
sYesLzpgjNzmtRar1VTLscNKIwaMOsKvZ5YiyqcPkjgTjD/UY20w+fE2Iz9orINa/4d+cHHIicbc
1gUabRUwoczF08+6skHNFfpFwlKmZxQRi5PEamhhFa5L50Gri0r25UqxKEYU53+j72gOEYJ3IrCP
P9khZ0LQAphPJfWmzVOtZuR/uc8cvbc8cN6T2aIBwF4+syX2xK+nKYKLjO2MFdEpyplRyr32s4SG
uRoBFQ7h3QUldztxbKuMOQ4HXd7aKLxC0omY7sMXXQ1Orf3BBo9RZ/KrVgCvTWeW7TnyN9LXdZ1X
h1yYs7CiAR7bO9bgFZm3NeHK0AaxS9ZcQEoTgyUCX/7E9+7NoQqZpNTstB03fIW8s8QQNLLo//JS
JcIpiTn6l4zR82wLql0vO65ZyR9JHB/u8m0zpGz7r48ZEvvwvHOuwYN69bcsDraykKM1s3a687LD
jW4PC0mYVeac8nY4tD2TUDDIVNcIgpxQk+4Sy5wkmW8LfE2BgorIwxh80Tv/wmDS2mwhZGmdyiD1
ZjqRhSg+t+soslmcaIlj/QLN/R/9vZN5v5BilcWCS+zatkun++3L0Sspvgk/xtaQtAfIoWXG7zgx
pAPbYYqEORt4v9769gfh+paztGhvYoxEUl/0pQ2qHUKibJNkt0WPZ8az4JknC2+pd1fghv5AQ7t8
Aan9NeZpK/hysx4WNeE2evTdnZe4VnHgldHEiQjhvGv5w0bv9UPuwK61UjmYgiiqm3oo5Fgp31U9
90jAYPgmLtGuDyjM9FEx5yL1K/eoaUYpCQXSwEgP9SXWVdJ6APDvZgizRErsUAmm3Dg0dWnqC5JM
NAV98PcNmiTrvsykpcfbVxhO6LEzaGCQotJcHQ6g1DBCSBJXRaHuU9RsZymgKvIcVtOC0JxnJUWD
y+bV2gVfXm64R+QLQ3evOrK4cjnIOvXIZy3ieiSgRdHuIqA4Qpl10OguEXV0gcq8I1Nvo0OZLuaw
e0fW4LMl4rHhjQv6KfdtILKv6cqVo6PbKhxFYizK0yE28yxJ5e4i3BvXv+kX0I9d/0/tzsNYTLxv
47Gc0RU1ytIIKkE7ZB6D3rOcvrcGGX26F8ve0orGVCEc4DlBG3tZpy4CGS49uHXa40Yent+wrhDf
g0nHGAQM3LAZ2J29/oIXYk3il2GGeBXMNgLHBHMMdjSPs5PCgWRfRqWJF6htWVq62XRCglp8mJ5u
vb1KpKYJF/Edn1OJPqkrbUnfi/kEPo9bIxe6GQZDGSwgZgDh60H7QUk8nrkPmmCsB5UyDDFdtbeg
m91wo1EOx/8MyQzBU3aQsJv711izGlmAIofcLhUF1uWpt92/Kn+4a4wGTZMc3S23qzxvW4YqprjF
6DSn0eX3Bx+ZgLF7fJJZFJqBKvl6oU6M6X6HJWEkrf0uzrbVkKgzI2XdcNCK+gg6G/Iky5CDMRNM
a1Pb2Kxe3kp9u2fq0sbZQYbKzCIuJSW5+PQECWNE91ATNZ2aL96Yed/R8Bl4b2mbhTRRnci/ETHQ
QGRS+FjlEOmz8qgbSGy7n2NKfwBeFOE2DfQQKQcnt20XHtWYS45KzHNOb3m0VaA8tBI79IinfFk4
JJQ2b0Rh3OrFmGw7u9OIdfbqfDq83KLlwsuLR/Tzr0dY+vPLe79t63JjBxc6bCYA4XFuV8ZOFy4B
Vo5AC4ELn+VR+hHv38fe1vBi33sE2/tC6Di6XDwkWyxJS0nvNiAetq8geXIRIVdaX7fq3lSXI47H
vxNpCXcV5DywKPX9JYOuWfi0QkpPh0PDnarn46IQ556twQvKmWafVa41dXDn7mCN5gNexVWXOnE+
980HcbsSRhPg7pedNVLkddDxBGJP+dHVTF8q7VgJiglWLk+DhuRO3kcIL6EtOuUyKyDODe/vLZFg
aFNQhUGHSx6CayvGBVQnATV2gy/Ifog8oMgj43k85riiApIlGAJbyKDlwfeO7gm7gvXRSYURImcc
TCog4MRd0MGmnJBFwU9kc1gtKW7GisFtH9R6TL7HEB+cykPVy3oAKKIorAffToLx1mXFFBGMoTjt
5e4ql/iPfPlN/U4NQKf3aQ05YF0zjEyaYriFCIyKBbnOaUoISUOzDFU5vtlnrtXhD1N+RfaSXN6p
nmuZTX/i9EmBAFPVYrKcaEsq2zBezxBgHrSnJDQGCBN6Rt/CoaXHB3rzGaEp92dEUAnd9mJTvDBk
LuecJkhIg/+qMZ55iqZnBESyu4nI9vlFnNTEphek0lhG78tHPcoQJ1nxJsLOaj6gkCuL9TRCzS5H
pWaTwjE401+87DEpI8Z26KTMFw+5MShiEF3okYz8kPqWkKT32nBeKMIkfxi1+93gT+qzKmFPAn2Z
nMipccLfrFyWCNyuYrfqkYF8hGp7dMMLHGL5jMLzjgpuSelMv7TlPLPHTyt1oGuTm7UmEsGDIvlo
Wp7Oq/YmwQi2Iv0bvVweIeSr93GuuTJrLF6+b4mG/2n5ckb89S1R/8K0gxN775Ka1CLSyizzcflC
7ozaISPc70lBDk68LOnPxfaa65BsTybhuCVVYR97mIsoeGKdEn8m4+Brs1KgrpsBBCC+8QvBx4+H
LlCia40sYOdPGzXDM1dztQtpM6BRMzcTaMGAnpOpdFLaai3/U6GIb54jGw3FvgktzDtYver3R1kD
Ar1EI0cMTW6Dp0tKA5ihpDL1FhxtxgkulIyTDa0tMDxgsuOKSJA9gLJdwG9yv86UGR3P43WoWA+V
9QxKXscrJsp0Nsp2cihC3R2lrDKMxxuDhvGODX3C+7cRy9cBR8EBiRWK0rNgqAnfJ4l/F4bo0xat
sGD9qce5nmZaDFz7TzMUD20PgXqF2CjkRiUxc/gXt3EMi8pnfcslQqj7JIpVmNbJ6IlpYtIUIvR9
n2rr4vW0tQ6rkdwI/EXUkIy3JShiYfDjV8PpFIaZTTGSs6CCHG3YQWsIRaMwiaiSQsH930DS3GqR
HXSGTWOAOYeZe2hrs5KlWXVXUAfkzbCOP4I+rv/W0NO0cgtcjZZn25FyYKLab+1WCdhH0SlZw9hU
AfiAlTIm6yHH3xC7CmJ22EbAY5ZQ/pMApFaCWs0XxZJi952a3h+5L2EaKsoqHN/7p2VqT4lA3gnn
vaI86q78xZUpvh6tZbBI3g1angTR5cHjo5MYV1W6rEEGvO/x6SjQcHgMHT5Kmn34jiogdpoC7MYP
AS7RVRAm0Q3kbu+wtziYMXd2kcwu1tXBtloNBTX668i6RtGaR41Odm01X82TtiNvVsmz+XQKr5M8
Bwnj7KusDPOa9s+aYqLhmjw/BUbR0rSQ7hVZAiLCxBGZ6tTVgUMDIXY9oDeVbx5WLpSb3DnGesvS
wn2rcp5ZLPLzf++270sWH7FC3u1biAxjiHXUVLxR7+UL4Wmr4Db3xNCQ6q+KalhPz6mGfHi4/BEz
oMe4j8QoT2L1HVnoi9LNXv9rArOMAFL0JhP5fcmlsVnE1b/RpVBIe0bMf7/IADI2KRdZz5KzP1nA
d6/ZntW34GQ3kmeO5Ru3b5QAqpxZTdt0DJMy9QQNH1aTuPJnQDNzG7tmowIC79f8sQtl63vyNDiE
xDa1kBs0whgvIMZkw7NHfLTLooxv68BsQ67Iy/yj9uzjK+yFLsMliWozYEMHJt4drIKSHSyzyrVh
IocGfi3vK15r/orRK7aJJcXYmbHQWDAt33chaKs7XeFbc+wFi7RoJ+QWGqQA+z01uxRokFt96Mbi
/v77RB4qbq46B9KeiEsedeUU18IMhU6dwYSdmyUDwEv78EDZrF1o6EM7ka2bU8s5iFTyIMESGeri
HdOmyQeMINW/d0tdZrsB3mTnGTWW+JMbSPGlnHyCo5XHQHspJp1afpZd+un5b5C2pjNicmVrCpg6
6JGfEhZ5DZ/ZdyOzdSkUZfj71jmNXK3PPMvRxPL6Zf9OQG42SKG9mATzbF36iRpwZy/x9W7pFN/Y
BafkAlxGC1KD8S9h0aE8FQL8mEA4YwwSNFcKRrbPdWdDHgE0KFcvfsbBR1xi+GKJAS8JabYTB3uN
RwNRwQqLbXDhfpiwUVAeegf0kAMI2J1ErIX+7pQbjb4pHaE2NgRCM2puiz5SiaqIZsF+7dSyb3ai
OdwWqWGrnEOkQ2kXSja5zzwjl/JDqk9Kkz3xYMwns6E1w81dw+FSJfmujc9eaXcXLoJd5zpwuBnM
4uKe0J0GstRPHVVUZrRoWwLL4UxM7mTa10ivN8W8KYbUEWMnsbtIiqjzdpONzAkqOZ4aFmbR3RVJ
p/2LECODdJzArYMl2XVBrURKDxEoQWFpbGGpmYtnqZ2odnRmj5n5wdHwd1HdfwQNyAJrQtjGUdEN
nNLyWxTyv7bkwNCPZf/p+ahhQdlreeGtzhLpABeUtxpVcR/aFvQGtJtuqMp2T80JCjsMrOWJygbO
TEkz/7F2yy1qGyHvxTGTUn8d9wIBsQQfj6ZS/WjXjyVab6TC4m+9JwczLDuTunNv/NMUp5jfCkcA
iFLw11uOdFSZI23MQnYD1mdNq9H0AC2aZ/HYeFsKeb+9VeUB32DJeYG31adzbu6GjRtRqiLy5TLe
g1MIVxN7NCvu48f0ukyXRiZgcrezDgPXr3Yeit6gT2Shg5ywQA8LPNlu7SejpHaf7bFVOh6p6UhL
l16H2BSky4F+W4sHeC7Y9Ui5j5vguRrOkpDe/OYMTFF5oNLsWb+1SUHmRmfdB7riVjH05vdk0pOj
7P1gDxQnZAwbIkPwaFsSEtuITDGJuL2RzPCJ66aPaDUGrOGl+CAdEqFPuouD5fnyeduDBDQI2MwW
WOAZy0S745HcFw1jx/+9azAGyPCzq7d0Tr7W0rMDCJWG6Wpjz78zGjMmHZh2d4vaepNwlJB1OQZ5
qD+K92rVlN3O/goAWgRTTnnG9uk1n9YqCzJmoyAtDs/7hDmrevGY7poVEzJ+WsB7tVm4QKHlVQR3
kMuad1VteL3VnjNVt43+4JduRz2WW8chKCocF36N7mSSxN2TeK35f6/PsPxT8d/bnt64cQw1s/vU
l3GytdiFnROjbKvT95WGW18t8KvhtKjwxSphHyTVJZy6bk8E5RsMeYHEQCyH583oIY2uidFzjRSb
tErbEWxB8OVeLHFLM3OgaS50UUJLFwx3nvipBPQSksgN0ZHAzlsFLNG6q2+xnuE2qTXRUcGOJFxq
uBKMkRvEIcnwtwj4EKeDTXKqXTVd47KbYVypi6q463FkoAUapAkP+7cJZvAYGcJupJdIct83MfOY
m6tX5COVOg/vtvn0p2EBgvikZnlMtUvBHq/PkD4HiHzgFIVXfBTIH8UhBDLubsfD2tKrI/bp/wHx
wV0ipD2GxrxBGuo+nRwmBdVqraLZr7nDdd3hFwsoOfQG0xAcRC+E/SSDyb2yHE/vrhg3Q2Mg/GKg
noVB4CHn3uimg9wd64nCjbdM4kuhTlxbJrsop/2IrT8r7hDJiguRAhHzwA4zQqoeeuWitaNCLmoA
XOgFg4fnAUMo3KvN44n95C3iJZcmm6o0qTZwe5tp4F+4rUUgC8hwcLYwB43kbfM3T7pVKm/TjEbt
DbB1Y7bYcqAfcUcrqDcDJl9Wken4cepqRQ73XPN2EcqRChmtYrUJ0694807yYUxO4I7OfM1g3F3o
t0wRezwpae8YzPKGIyAVfCqEhTSEMBoqgI/ENr1uIhCI3NgH1XgV2vpXVFQTZ/BOrSgwBNLsyptB
Lu+vH4QsWLxFYFoAA2OGhZVo1zFWqblL/KLTimQhJO6MqE/wW8EFv84NQgLF64/mgaXtaawjsJKz
UEZrJSTROBftRvY9wC8X+OVUE0cGeww/Ew0MAPVRCdyEHTYke+uE90Pzmb5NYkIxwrBDny3ScusS
rTo4wZ0xea8hzamh0qZ09PZyV/guhg5QqXIYp7Ou2CpIqCUpdFWLZf3nlOhcaHGDNh56TXSdVK3B
Vqibyh+2WosILtAKNZB8PfVAN3EpEPzoes9hcEMZZxwi2rYKMJ/bmT4czPHfRSMt7jCCTX0g18Dc
b2CZ68c9dWxE82FYGoVkDFAQe4xFSGrauRzYGIXn3HM1dLH4f5Qujz5KRf0ATFv+Jqq6ZEFdXtiI
0VKyEyFvA7cLMVcmQ/OrIcSykrIUTvPHptX+PvesqZar+2+svB551jwSJ09t2JdZH92LRDsAZvIe
WDzZ8l6AnfS8HARsC/dDvVUV2AV9GVvtlwnIYJYiTiwbDWHL7iDoJCdjPQ0tn9xhfyXEgRABkrLz
WjwTdr6TfGfa8TSjUEwO7Gwl04UPkMJhNkG4G0+s/D9nQ90YQdEEqOtLEgajkQlQFOD2CILujCqm
SHdMwzJsAvVJUwjmKIH7Zn2s6Kzx1zOfUPaCJmQRO6n33x1jIToGxuqKBq2b2ktH4dYAbbm4GiFq
2ZThcIAv8lmf+e97Gm07EfNcr97W255NTqVOX2SkpYF1d2CFiTfC1+GLkee1uBir3nWbhm5UcPBK
S/uHRC+hvsjza7Ze5CaoVgpE1WIRJIbVvzP+tmFrl1FqBVez9xNmsJK8I+PyLJe6HBYHdMDa7bSi
FHkQtDso3R3FMv3yDWaRsN+NWV76VbeB2PMGUB4HoZ4igNQzkKPa9YYptXwHmtUcfF5gtdFPPrge
ARPE8AY//Ia0ObZRd7ioiQBH/e5JXb2q+e3eGu4fp37Ims7c5KJgES0lqY4RMM1f/O7UqEYTafXv
sPupwU8b3nJ7ZNdc7QsFezRVmxYDX+QbufJPbsz/C426K/CdKmksZLL4I4xaspYvP9QjS/r/z4Xg
A7ejj/XEoeDGrTiwy9cHpn9d2B2blax0GB37ugp5pkPUs+ppn2wX1ScEzzPxSbD8g4tMhiIryNwY
dsXC5SIZzzQHUrZKoDIeVDflWOQBJOhIZyRYYvbHJSsmTPRaRZ52b5GlY2n7wUwE9/f1HLISPP7p
KJdW3puoAhYH75f6h5HcgKPfDfylKxVwX9KdQf4BpHiYFXoByZvVmZwxYTYAdZd+l7/4MbrdaF8U
jE1WYTQC2NUu55TZzFnQxSI+pd2Yh/ixLNZ/rjpqJCtt38dcucnyIGzLjwNAE01LxL8CX7abx3zx
kSJbxbK0hOKKwpAnLdfq667wLgkgw/zQxkw/3dcw+lHLnc4CUZl+TBusHdDJ6oKHyQSbJ2bgenL6
nJsDdW4akZOXmiqYf6vRhbfP8hhlwW0WY3oq9ZRhyliboVfA/GwjUNEfbXKKkS9p5eK0abll4lKB
mpNq0mWkA4UDd7mCNeeNVqFuPQq9VD3wBCL6Cuf8eb0j6JHCcSiPgKZh1WQXHDikp5KmV9HzR3Ud
j3wO617FptBGL/H/fdlF5+WIzP95EKiAc910GmVHWbCIaSzmQHRTlkds3kJIDqtWT6iwWc52qPwh
JvMtTAYuIK13/PCwARW69RwasC4LEaF2BsYiyHTZzsWbpgNT3aMCHCKZ+izdy8su4bB7+faKdBOa
TeCX/kPyvq2dpODr2jIsUNNqB+YLPYC8IRRVFx1VyEJDTFBLEsggrcZknlJGhECPFYj4ipNNBOWJ
wSPMALDMaE10N8gLVeWO3wLMX6aDFx9xI0gTVImC+COvLIt8rE/3PcTzjxw0AwfwCdctPTK8f8Ge
Gp2Qh1sLXMK28zBY8daQcZ5vffrMQvgswlKOX+4l1wk4boOlxyWrCe4bpF02TdqZzYGzYIkyU1Dk
xi0TQkSlonGgNGALiPKHhfMquiMWTe8Z0s3eNkA7cTZ3iYTPqizqj6s7fugysQcOigZGG/Ki4pew
VM6XLuxQ0SR4XkoKKbo5Obk7FZH0WO9cKWkM+U/Iw/14czjKqJvAqWE7mK/ZoKKVVrw++adbnNUP
mGeppU7Rlsu34GtwlNNO+F7tmk7mWcEfZMA7iNHR6jM+s0L+CKP7XqZrQlUJc9INAuYVD2yhWI1M
0aDqcP3UWI1+f5Qw2O48a7+mr9LSxqtxVwgqCzkhlMp5aO3YDl0H7taSzfSpxgAnVFSdj/S5MZsJ
WBCftPgEmn9rLuDBa8IJgIFhHTW8TDyRMBh24faOnt7qKJt/0jGxkghog5tC4+1ieXwP8CqVCv3/
H9/zMrZlu7dEDl6jH7XQKWjdxPDOWmgpIcTL0L/PQOwntncKnVKt40nrykiaoN4JtSpXbH9gKk9H
A5/VJ1GtRkvLOsZ0CeV6Ar6evBkgo1Y73em2c9bvXsQ98DOMDR19LYFU8MIVutDKynJ/BPz6O51q
x7NfWMeleQk6P4aJwdRDGczRZYXCyBVSg5OD2V07/elUKpe9tB4TP8LqtkVnnqfjq81udT+rjaPv
W8cSjYRwNF4NnSFGiZ9huh7tjKohEc+bcW2G0cIhaaX3G7p79+Wl0pbE2fSkaRCwe2PL7l7Z39VN
YRKk6kh32UjWWXTZ3QR/LEgptkOGeLJ8HotfGbjK3u5t0lM5sZWu0LUMArOeYcidBOUfOOPTbEzp
9E+pb6wv2sKZV2Ff41dIt24e6sdyTXnQ7AdGj7lB2gCdb4UnzblrI2N18kJf8L33x6rCbXiH1+Fq
dbCj3uUldwTEIkLijGygKXEycWE+JqDN5Ox20uHoTUu+VsPC2Cu1YeiTlDpYXXx3EoWWmsoMN9bg
CdrT5ue4GPMK4VXd4z9Jn+8XvgfEYjvRRtPYKG9PuDA6mPoAOg7157DVxJVJw2w3xJ2JBZ7qEuqg
p5sH59SbZ3+sxajnPJpK2u/NLLnGij8tdWnCh60fdqWWNn1Pk93ab3+75w0ggy8gUHtvcV65hMxR
P9kdWSmm7EBFI0+4CLWB4M0vz09PSP/Wbem04sYd+HYQ/MDZujAxnJHzWGVn7gkmUA6e+y4EXhE3
xzcFIjc62Culu5sseqiWVWjOchphY0EWVv7C30Cc/5pV2tg0gjTmyIstNTW2uP9E5ZlEw3N5gv8G
CJVdlTdbGzCq1kyfVR3gnWMpF76OxTHuuqjzYXybzkKbg+QK8lLg7GieCElp/i96y6as/Tb6R9Cm
Zme5DAzZlNQZEbbG2fttBpHlLhUWZk3gMWDijC3wfrAKwmuGCK/tK/wLA8FteyBNFp/JGFGWSePO
xkvI0ePTLHNa+ryOi3RMMR1SHUklbPBiprEJegrDMJObY1O4xXYX1kOWH01iFSnso5f6vzJbfWAg
HeSS4u8ps+EdrDn6fSSEBtP3Lh7q6jCgjlEArllS4Bg416qBuX1gX4xddSq8AuEJ9NNyk6U4/1T/
9q2zS+7Yyy0lFUHxK0ttJENJAPqzydBwpoZNrOYn/YzYJJ+kCCP0LbdTTk2UUmbkEr7Q5rNgBRvC
OtH6Sx4lPmTSwd9PwmGQqHMlzKOrrb2sehDsJq2Lml9YBU2rFQ6cniJl7/Olmm0XVyY0vD944M5d
y5omI/t4ckTCeAkK/OUSOGFPBeoL4WOq8Pfpek0ujQEQxzviaYhi0wTLDnmWFGhmOEoDBQayMVGr
P4EdWhuyKvxmePo5aQpBnjBi4BryDxWGp0mZPkFRIIy1vCzCco+2HouDe9JSHO5vejIj0t0LNtuA
PSKCf8YbcDjGDtuVH4P5Sr58G7bab9FP7shxX2us5oImsdr3vyO+p14pDeE8VUml1PAxw7TPFBbU
3oHpHld+ng4ITBPRhFh8UkIikhKTmFxKoxizCWYOAwRUwo0E+T8UWWzEgOJDu+Qsp3wQEbgG9wLD
o6BnKZwgLNPHvXpu2oMH0dop+VnJvlQ4lW+a8ErNBbq/vOaMOnkzOGjjw7JC/XgoXzZ4wmUbhOSL
e1VwFIp//tM92x3EGePy6MM+KL3QDsN8Vs9GRFepoN8i0uoMAV2qv1Gnif+5cYQ13Y6dGxUgISvL
b1UyYcaDuTmhUifPLFsnHm30bTnog9lMGXNfCIFXvuzULWpa6+qoV7XmZTyQfPrNDnEMpX+nIdOd
9/2O9vj+5GQSLhgxFF661nebgNLzHGSWOwz3jQ0naprP5kVQVokZFc40R5/jUldMow5xqwFnRrzC
Ma6RpQXoeUJnp5DLt8U78oDzBJrup1b8azyu9axvdwSF7FY5N2GOx8nA1YFJpq8kdSoC9tTHmO27
X1TJB6kpQ+Sm4dtAfLhKGQqzzSro8dVXI2ayskwsTT7JPEeWksV45gHW3pulTUjUwDZ7vK29sF9h
jQtVK+HHhb07eZtl086CVG5pfiIU/Kpt4BBNmH/TgTXmQFxXBOIZyBvpReVHHg4/5J5qh6i0XBqT
qeESbZS0E29aizOJaVoiwmSLTOybEkU/cxsZv03fJKtZW4QE+QiTorY2G3dFgAEeWmHg+AwzX5xm
Uqkm83+iCQhj0u9DFSeTZTIVIzn2fcNw3ifFCoNDq9HU/e200hiTBCcZaESARRaQ+pF1KZJ82e3i
uUI637xhRpPSvgktuIhRvoX1MLY1Xe7XvsW/Baf5zQ5jmfh8gXI0WIKic/h9lvC43HHZn8FCLFUJ
lhlFH2+uuvM1fs+Ld6u1xtfqDSL1gL3bug7Hv8Fev7NQSB3LJluZkmLS15GJMoNLpylLJThysFA6
WjLzL/ODqL91kmeXkFnj7X+Vt50qoaIFns++9Gd0nIA2DGL7Ny5AWUxfMmpq0SEAz3QWXZ5y9C/l
gNytK6z7WtNLfIve7wqLsk+zWLxfbEj22+Dw0/2QrAZGXvtXIvjNGw7uF0WIERPSlwNFEBri78QQ
Gvargw9/xeF8nkcRppyg9ZdU/kAqjbh9EWHoOvdqPUJP1qSzqN7gETiZSvWOOWh5XFt4NOwbMcJK
ps1fApeQK8erG9qJ2G/PWkODSPqAe3vM+SaLXl5jrpVOcyLkTdj6F1ygc7DK5/5mKMJ/JfDJ2xkW
Dg8h9yrQATlquOhTKjzlWHw06kfYrqsGaAHwiCVjgeT1kC5oRVlxqjcW6YMbEGXfqv6+DA+cOm1Q
Gau60JRSf4CSLftD1vCFYGQqqJr9A3LxStEWifopt8s5zVWg+eAzzIy1WWco7GZILNBNWbhZa2yw
Vm7xySYRFSJwcl/BaCDk7PyS/x87zIKe8wVBXXSFwxNFsX11/zK5n88MIYCTcxq8abXybULR0cDT
Y2K72NvM3TzvcK2KEct/W6II/Ct4zWwn0gjFKJdize39emByz6krbNjC3DH0Lvorj9tMqjGTfJ6E
yN/XTXsun9OLNxIaq8A9ga0nMVVnyR2hnVw1Mf/KFAi0vzabv6aKRLmT7GdhL6MgvhaeXpY//FOS
Ue/j/VSXCUNe27aIq6Co45g3j8+mhTPU4TZ46f3fNiwsFNtCzoEubXUyREFpF6bok+ex9CLBuMYc
qqIm5s4+oiD3fAWGuSa3hkoSgPLwaGg0P/JNDyA0nt++8wDRt18lJct4Y20Zj0kaHeJ9peusX9Xj
oCkYrEIkITFgRby41BMb6qWJAyiC9dILhERgz7gCkXyBUC2Sc2+RrhlzgpZRgCtIWTHhthCKWb0B
UtW8j9g5LhjyE9tJHcP2eN7vNdyz6sXRnhz93pwCM3JLy30O4KhhFyvD/XCPXQCI08qIr7TbuoI2
OgZ6340pdW19USvS5nadtxkGpxIFrBUuZ04U6XuatwwOMVhSWbpxKUNbVS5WY6b5YBhouadOEZRw
JDsPLs56IOgU+GzrB1PQ84EFRipjTxwiscz9r/jQWAGyi46wUaoaBPob7eITeUAeNoRKreqvrDyl
4bfKU2X54eJpfT96PXkLnRH0UkYbPzdhOLT1QLz1l5JZ4ZCAxoYHxVTm4I+uuZcTEhh7S4jH8QzO
8PKvlwxTT/c9kUqzKiYYblwkaqhTOOQBJpyeK847+pgwBqJ86asIH4AR4mWyBVp/YODvpIJEuy3c
+3cZXow6aXwwNQeRpfHt+4Q7ZxHMKigwdpi8+kQ1s6XQgzuZZAuJEP3t0eUhtkmx4ZXmjnrijCeb
c/hLI6WEjsjz5mjIGpVyaXCISo13TbLP6e4Uy3QUZBhnr2mFpap7NBH3ATVF8ozwIOvLimoigwaB
z3ryWRDv1Wf4Jz7kHpAshsQDh0J2HX83bYG6nFsuJgTze9esW4OMSCVPn3zvbQFn8xZMoha5UOjP
DhfkOUmCgIDFjwDsgAYF4ytbURQuSIxbFD785bbsTcoiP2fI1Zz8AJwObV51iiGtYCD2U8hH8NaI
GetL8zmlx8TAT2fZ0JnNuNMFwrTJ7V0SQivKyZl9Y5RvkJVUyKEeYFzfpgTGmky6EXsUVUSR1bTv
ER5HYdl+SqWNa2jUkS9A6ebjQ73ft2wZ+F1EyHtOdkuXK3QCqF7PdKim7pC8rit1fBU02BzxrZbs
+aZhCk9lcwCQ5V08h625nsgIlp1jefIaj2ZhzzVJsmq4Jz9CV2/WFx9Jo1bIF6fUEZSGaHAquO5t
1euanfiWYBoH4iIGV04KXzMwK+BoMyp3rViaGCLwi1VXf9tCM+fwN2zNBPwH0TlWyaZzRAjWokkU
UmIZEN6ZFK7Me+dlX4nN3/zZAmrAirEGf3WydxODMv6tOR6PrrPlk0NYu5+u2ViogYkzBxsHD/H6
ltTULEg065kpenPgRyVZCugcgE+KgjE2XADbnOGBJwwK6Lvww/QJswUcadzp+bw/7kLnGwrie3JU
ls0AsXoYhK9DeDcd7SlEcTrK/0GF/Caw/TTg9fsVjXrcvZdk/NJeXraSESEA8ZDLMBYN/+VbpdQV
QtsfJQG/xhmHv3XgpJPzAHc4vJoTkzuem58HuGGcHyI+hhAe9G+lRORAoBaqXmojl8y0CPtSuXuP
msWbRMUy8zqlqZqS/V/kP6BjJCnR5rY/aw4zWgaCKUhSksrJRqj27MW6IrpO3ftp9miooCNaqgVL
rgttarK3Iflr+d5KOb8O6JS3oKanR4BjMNMRVib8c5MTE9+tIr9DHrinECAbU2Dz5eRnZCxgNg2q
QZcE+oYHMlHUrzoork/t5mTdfOjV2ifmw4rmA47Hl5AmlwX+bhRSEVCArFjnEXX9op6Sx+TaGykh
2k3kcKooZ8Crmfeg24mfOsHiwv1a1b0CBlMRBmgWSkEa16IKkuNx1OBQYhVIK/pVoGFAnyOxOg9X
BlWG5QNiiukByFRUTS3B1dh8mutni2kTpPymgXLoQM0dtQWcLZB/Ymzr5tBIn6s+suEc8yrZ8klD
4bDR65oVy0Q2mzhQKZOblRCnKRkjrEpyNxbiLYwzruVC5nf1wh+dJ2EObS439LbE3PwWx02Yj2nF
wezQENm5+qdufJQbPpT6wXk0+99YwfdYZ1+kykc2J7fOx/71sojyjv10/NRKO9AFyAUdnDEEtXjm
JXFbFDL+ltInnh/ixG/4iuGe4W5jF93wOp25cLzqOInYJ1CRmS48R24GWIp2B4aDwg9LUUZngTQ/
O8f5cM3ElgRT5K6mBnI+tc4hRXKPzt837DaUJVi90i+VErQxXEvrupLkh0TXcWMCdBDY0yyDRB0N
0r6ChYYC7NHiDOtQyfBib2CqtsYhakV04rpUpQM82/sBzrh9WvhkBxCyUW16KimKAvKdX6CijGm4
qHmU4Ici+WtV+dAEjgNgL96Nd891ts0/ayrRP2npjlto8dU3oaw1pb7Q4+itedqNRUYqEQGSPEjl
orfYrqJu2it7XkutuyhiPRLAtJWHOwuz3eTymddqGYUqTG+o0poz4UnNJnu4uNV6zdrLbp/41Ave
r+oVuo5fCPBVbizV4V/4s0jhl5+X90xI2+tFXL7DTYlbgDyT0GBhHrEd7zkFM5Zxmwq5zN5AkNGw
W9DvKmo4WyVW7ocM21hr8VwwIEDOptspLirohGHpP+5xOhLYbEOyTi5kIB+vNov2D++C6vEaceEJ
lPkOxDwxgzxNkHoS/lqSUWWL8qkS/chgsjGC/tHda1lQvTBUGTbcxh4x3w3i2u8Fez2yvNVEA6aB
gR5cmHpGKFJJ1B/Vn8+be4wkFECdE+VV6lI19nVjyo2qAOW8qJbpXl8s5VzSsN989wcMGykUeIl+
1tldD4WopWLI+lgWcZbceGsx5I+KSA/OiFkazbIpV7n8x35ir8I2/pej8Zu+MxxoIqrwsFZKpU7E
dYu/W1BTyMDIr7xEtuDO0uXLfw5EcN9R1uMVljXXlUOj+35wvFgI3yxpGGqUmCSIherqeiglccqD
V7n8unKFu2+/vJcCIrnfInh3pqz+Kzp0qaUAHIQxlXAsJHObbJW4PVJsWWnZ8/5mlSNLGFloD84F
R/cNX60oeaINgGsaVURuLIv7V1wP4n/ALI/ZRCT3GjYLoxNmjpXMLWuPSsM6xO1uxg+rT5k0F5On
wKfLthlZjz0mOwAqCd+jz3Qxp1aGjfjXu3To2FGFM5xH+k3ViuzOXqAy7FEaxJYjQBVMoMa92T1J
LIKApm/v58KKnpfV6WWHkJcG1VG07RO2xs4i78P+O0pdQxU+/VCqNv9NqRqGaYOWjZnb+XyQd6TS
lzSD1qGVuSPvXQ0EGdymXZCUNjfST2rtPwjgIB0zfWhtsCu6b4eGHbvTfjBuJUwWgcbI5xYrS1ex
WRYnfvSvOyQlB0luHYO2BR2HhbYsi0dS5KtawGW1JvDOufwaNIYvRkn3F3KdlyRkrtfCapjoUSUC
HQfnwXgoeV/RlYmltJ0aqN0RIPG+MlaJJVOsVJq4CnwffEyNSKwh9uy4Ka8WzEygud2F3JEiV/sA
aUvkt5eU9CFVH5ruvTO5tmZH7gSgugKFUYNJOVrne1UgIWnxSB/e2M1CrHH3D7UUageLRmxRRza3
I7j9FgCxi3nxFjX/Q8RcsezYQeXpnyAeIb74z3UAWN2rYxOJi+omZoS7HuX2f36emofK9hF2Y7Lx
ySFLleJYyPkORsfhT49kQZVqPfZrIOShsgNScDfiFtmqy7CJ4j8PxJb5U1Y0fdZY25QEL1qfBwCW
jP/EzxTsDEvVDN+8v2gudAS6SFOEA6CnAOyWP62jEeWNAYXnI/oV4CefhHj/AX4embzSFdKxy+O4
PPydyOwkZW3cBsb4XloFL0E5CQhOuJg4LsyukdEDGY5Af19SK+zV85v7cTqzFDagFV1Giz2KBi5f
vFGbsj/Vrd631SDoPs9nDz7uqT6pO1Um4waIEDCEES5/R0jXseSQfFk6vdgM6HiK4dP/q9Jyudmn
cYpVy/DOGzg474rnZw/yBlsZYf5yFv1JelvGyr53pLtQFKdEPfMzAMn7/z/bqkT9koefha6+9sTM
HqcNbTyeVuI3zpziXi7EuzgLd6FMZk5S8pAR/PqxVtZf81uJfbYiCcHpbPyFy2VEU/bJ8j5iFqYq
Iwfa3ipCK1p2mRqz0K9kO0tCxDASicf35tw75mhaiW+piv5ZTOCopZmwhBrgKpVX3hyTeG/KQZ2y
qHbFJWlAqkjGb44VQBkfW5MvHf4y2AiQGjX93o7K1KWiF2D6avwc8RKMdb6s0GtDPrVzQzYjHHFs
LHO2SoP67qnLu1mz92jmJcwKNts4D74nfRkk+JBtML+ni0OlZEaKGyLJ6C3zQsrBSpaN5gagkxcm
+ZownwXX+nXmF5H6GMDGMBk5AfQaapvhlMWX7kuv7QTP+m+00DmJQtisNwNYnWBwcErMEKD21aP5
XQ1eeZsMagDBQ/FI9C84/KN8+smGRM3/y2jzLjEC3JNh/Zm3mYJh7Iy8VY/L/dvdbzfyMCGNF4ig
Cmf/vV1ohjPwz6NmV9kZ2OV8X2S5XDBLpoC2d0NddtXlCSvy/euDVTu29lCtNyrBKJgRO+7si6i3
FdsnK/hQ7LYEYoxr3rtypDkNEc2/XmFYzIqSXs4zQUCSVWKdxvbKfZ2CucuiXtfpq7mOisOe3eZ1
WFODvzzxdwmoh5v5JjfCskL13HgN2nP7fsdgDsuehSGTD+gLgnxo0dMBRPR1xc370Ok0360i5KdZ
wBx/C16nSknCAT49JfKOlErbgcIx+juSOzFDhH0h+KlF0G4tHfv4AjdMCjhkqKhKi3adIQZix8Iv
BxXATa4u4ohyceu1n3h+jVYvSf6tv9DojNLn7R5cu8fV4eFIT4udYwMBcv+LhGP/GKk/KRfPEqtv
2YGzzpoUZsSAu9WPSGW7omt89iBwLjUILeGOkXTVDgCx2CDJ/xX+hNoqA5hOvwRVwDIEB8XRuP06
7B+wBN66HiQQGUPuchLoMzdyVAA77x/ehc4JvatjaXru0ttWqO2JaAF5bk0ctgBC2awNWXXhJvw3
rc7SwhlAwCWGq44dN6/ZK/HmUJEY69S4xi56m8x/ysGNy8UBAmW/GOAthF0Jj7DC4xCdfAVp+55E
c6/RbyPzaLfjLDeKDLFs9iBzp+I6O28vYr/4pnisZf23zghcq8zq/OxpDTwWIpVTxj4rS1bfqLiR
DPcBZZMo0y4GIpZWFP/ieb2wUHT06iHVDrq8jZ4TzxOd4vXjT0YMf7mcDE/qNmXzxl2pDwd/ybCT
yK4cZHdYAeT6snLJPJgRndlG3aCf81YPWY0JZ5TTVHcmNpxq8JWx7EwETEGwc+UkmT2oY0g3pXjO
pmhfJMA7YMjjT9cafvqq0CKs+Mz7ZjQoTBs/z5EjKOQEB6RR7H01qJk5H/BK6qNFNhVx7pu8aEWl
i9x4SFl72JrIhPYX2+w4DwbGS3ALNLflYny4MsnQ5fe7VNb8CTASvzancGF8oGynyVxHO2d+V1t6
yfnpM1iqPDsul/hljNjtt2TaGsm3Rr1vVP8M1sS646/o3H75awzqfT1A1Ca+T3rIx+hIAWAYt49W
R4XJDeEd0+F//wxDZXBZej78LQQqbYLAl7VzuWHkqBC5LK9L5IMT8G+lbWlYCgGnl1jQ5SxhYLbL
lC1Zo6lzgdsC9i7NLy3AUyS/lsQk06LIkmh1bEGGSEq1R81C35pXyIjQvWvz007zftcNLDeJFEZB
uTHQzejJrmtGB6sZA8xamez66lPxkpvshJBnC2ODMYq62O0yFN++R9jzZARop17qgjpsQJ57oMQb
/lLNCfU7sTCXkgE/S8hK/C90bjEWdUqLLBbMtfizJJ6c+SOMakZdcqIkfIyyTXRTILkSClexi6cF
tj4QX1ZEuig6fFCWrcihPEIPfwIXYBk9on66KM34S/gC6W3tzwltDAWxKX/tymcc8ln7+ExW2wjG
ykVG0eTj+pKyCIsNXmNE+XMkGUqwkk2uRZEjUnM32B39+l2ieB18t384n+a2j0kN5OEDPKLMVfjB
EImn0GdmQQLo0SnfGBnQKNMSwrsePm7voyqRT1rREL80g05yUDKO7cMYFtKstZ8p0NhLiXiu7P1u
MyxXBdFv/UFHEDk+TcVmXBhKiTJfSXw+9sUaLt9/CJDH5Fz0hAhXFXD3jsgZJFUOhNzM4DXDJAX0
ch+9CrQPNXLW2trVQZElrpj5zNpaCTuJVf5Lx2Po7ad6oInPcokKJXrKj7WfdOzumMcYMlSZQQPN
ucAfZXu0i9IuD+X8iv8s6V1jo+fT6OWr3AjZxncD6Mb67rccesBx3ACyukWm5On9kj3sC+zK/Hgn
RSMJi3mJWxuaue0KNrMNGTO/ClP5eMSZDXGeoAp9GlrsBlUtPU0iaplxAQfRR4dTiOYQae6LbQ8k
Xw8TCGfuGzLtg9o/nqBg8s41FH6fq5qZBE/ApiC+YVfAitlpeB0odXInLK5IXXSo14OG0h3WixYn
5ggmxn5e7shciQuCEUFDaj/BFwt4Svx6xiuJmDKtyU3GTmWpss8pZT4Y52VK+/DXT1OOsRtub2Ze
GAGaPoHwcOOcd430+SrJVqm+YL7BoHaP9nafLIKpAHk/dKUlM/bn+bFBjnKwVWTITqGS01/Gjxnn
uFiuo+lPHKLvBkNZE1a74Ldo8S31AjK2AZSYcXdMGQcp3CQtw67ArtlacW4lQc1dr5mg3jo/ByoO
1IwKiByjI7GDkudFGLvYbR4NkBJ+aCekAhfzx8rN0xLNjB0UniAMhD6p976i4GW7xBv6NjjrDA2T
sPzcsIWynjSMMq1Ydt5iOwkp1iXujD+fw3KmQAbzLJEWrdov0QRYM90yU6WaEax0B3GiwrkxPxXl
73vhEedk4PR4oHH65xvzx8CDiHJZUqQWUFR7jBjHq9/M3W7KyjWxaQCaN9AAjkHxOD1a204d2RwZ
/t9FOxbcOhPFdJWI/ZeQa2kLhhrXLhKAY/jWI+WclHzb2bUyntJI7blqHhQ8p5LoL+prf2IYkEfk
+W85VTS8/2ZBnWKbxBoxiwSXxZ+rPlbG2AGUR+kVowTDzM7hrsETbd4L4FrUpy8nMznSL58PqHn9
PFRsX2jN05JcTSbBcDRf0pFm5v5pUi96IuKpJ7Iam0FHXDGRcyhpywxjpwsupbV6Guw1QqHCuLF1
w0+fbQAjTZg6tgQGcn1UMHRRFxTfu5rIdy3JFQCULt9cDzxSbuIR+do68N7TThRb6Eokm+lWbEe0
heM/7MO/BVOyPg1lonLP0UEBzZbwj45uFb86NmSwYwuGkChl/wB8bZKU8hnTtm3+Mjxgm81aMcM8
a/KtOEJXOMCH2UnXH7i2Fo6x8mOK/Zjp6EJ1jqkfi8oBAiVxkPKY00Koh5qhX0wezMkQ+p1gLp9x
bYmddsNKv81OQvp1xcrpUmEcblBbZLhYMLyIraU4pcZdCr/KRrSY82tZdSZ9MVMPSa96EpJOE1Aj
EVCAeU4oZQzBL5+UCOxF4puL80+v1+glCqFCiU9cGoDiSbR08LSlQrt3KdyEaBwK/Efbsiib0+NM
ZU0rAUqxodLuI6esBkAWfCVfz+ms7eJwFjz+OKoF9JY3raRn5PEl//9zlzwju9YpmySSIsmHoUGA
bSAba7GDen+Ruv2Fw3ZvU6ev+3eqFpEceRi4OfIXwSwoX2qlDnklnYflUHrHlVkuvN4D+rtXyxzl
SJQbyhFVVvgM4CPb8zCks3rHztBKBxvXLpwMgVo8MZxYGEJxI8fQR8R3OTBu7QoJ6HdRt08BnOtt
MWFJUPlgMIlfJMSRVeDmmJNthCtLMyzYD+J3UzmUMqlpUGz/YxWp24D+E4aIESXKUNfV0FfGqgaY
BFdlFxSOrFJC7Ct5YQM9N3C1jnSIJbS1beXEwyfHrSh5ATmSabbL6NTywUOHwMpdinOCSIIUkg4D
TPcsvLSKSCiZAelISvzsJIjJx1a8l5/6IDkUFfkUmNH7yh+Q2MfKoVVQ+PZMHaTclh78UlnSgMih
t60JNGgNSKn/rb8p2o1ftniOXLrEzdFV2TJVZ5xtkUENlUZtc7EVs3U6wGLr8vwJ7ym80nQuBe37
1n2pBLVJoMPX2owjKpB+jxZmenhrlRmTnZHP+7zfFugMx7Ob2565oQbXBaOzYnTOOMm4rN/253lT
6YL0nbnycFvf3faGtxjWnALyVJpfiIdyPpEHnoqS8hayqkCFtq2JW7YiA2yVThawmnBn86IWcau/
gQQjKcBJtXhn0ixwI3IU4gaYbwkeBstu/k4WRbLKeXgxGPnfiF0LyXrEXMKBs7OwkLJxEqAqhDUc
rZheBnJzCh+SxIJv981a2C0nudUWGBm0vrsrELLQR6v4zeezVmtf0SiqQZdw+RPFb1SrqoQBsYIQ
MI897mWrgS7klMWk96D0UNk9I1ghD8wXLIH0S+Ly0Oxq5x3iqW0Xk+wgL1r5BTvQMdRoNAH2mY5j
WZCNyrjMT2QBglVYOzxmtwOoh115hrK5Gefmie3YBMEqLmjQNO9GEvg5Hf823qypzi/c7i6ciSdx
ya7f4mLg6YYgOGh7dREd5hqhOeYq0n0J6hC5t3OXVq2I9r71W7XdoFl4SAP/0MljH44UVCgm4sAo
fpvPCspLaa11E8zeh/O/xzN5zagzHnL3EpvXyXa8NVX5xmgNnpEdztQsBbG6oi/kbpMpY4Sq3LfC
KLEYs9ze2qrGAAT6MXrDG49RShxchZTu1zMnMMwD4ZQ3TuDVczByAgye+B/J/CCYnFscXCOmcrid
vszyKeMHqrDVO0DukI1keBxSq2plMjN7KOij7IDBvUYKjTeSBD2CnvIIRwQneUPe82GNWbchiUJf
uUmpaBEELl76ZL3sDOJN4KFGcKH2n67XU2l5BuhZCZsl5Ja2BLbaj7KpHehp3Io7XQ8mbmGi1q6N
fWKWtxD3f8g9NqZr1tElgIGsuS1g+ECFFr3ob1YJyFKp1G6dfHyuWbWUSfzQqRQzUnsOEzsvmeIq
Gu6qT7kAg/qVkuXMtxR0cMZRjiEAGRzfrOWmwrIWeyiS7Lb11IIEaEIz7jO1aJaYCiolahvoUYgn
r10VOku/SjaA0mjvO1jZ/0OaG+SGH76erfDHhNJL732e89WBqnenobNfIiPJzD+Y2J7+l8SN4YP6
l+rgGh/hV21vB4U8brLhqphwYgq+y4ghUUUZJlc53XQunKyzXWZ31EdKDjTzgGk/GB3Zc9Qb71At
yekQCqExsnQwEa6KgoPx8Vt7YCobO/wVm/CR13tghPdrVV2q0z2XabY5B3BvTEFVotBtqenUjEm/
ni/1SzoJUuSxHELTG4ZGGtv6ogZOBOTrBio7icbFzR462vjHRUdAmFl3lPr5c5qj+TUEThHDbYa0
cYfR8/Mvzgket8wGDzjCnla4ZujocTjon+twxOq4F8WagtJo2lEXpwTTrfVvnlDpH1bnR43KvuYs
HE3XaVaeAFClj+ubfSD9UNHxrCnrkrVaKAhbT1K1Z78LQDdpXs1ib3SDDJlGlc52HylOKxtgbVQ5
PAxZlqL2kd8AoDSnkiv7zRxwW5QRZv0Bfx6UxxHms0mDRGNPYSMRxFBY9uKPrAbmGnsqb3oV/AOh
ixEiLxUpTtY5j0TtEZoiZ99cX/QHvWA8Wj2fI273izloFr+mc+Acfn+0nr0ktML04QorkDMT/lHB
8KlGwEHrAJEkFCN6tsl+jPvhSKYTsekAvb23ijzOxN1Gv34P7Ms7sxid2MztdhfxjCNOa0SbLzRY
mkEDM1gTJZYZLUiNS0B1N8jIf1p53EcGedNQTX4PVwrZ2tkrriKRSrbwr+qoHpxiZ74wGy7WkuiQ
XYT2w1oILKTnzauuwVegoznEIk71l5r7YOY51ne104lWm44mamFL7CveFMen66op/yMXZgt/aYN9
DmHcHyScqjuh8uomAqnS5f5a/euDhNdbWQ14ibSSQ0Rt9wC4IIVRJtgXGnlbfn5vaCCAIPfO+Zcw
yal1XSO5Sgll97MvRgvl/r4Afsf/Ru20xTAeVcr09Y2INAm8Ue497U7nKj1fKdCpvMhOWDnMjC4T
VQmIIpB74NsrTy9QUC9HWfPRTId3v2wKMY4S51dR45kWOXk32bs4o3VlsarNLiqvzUBceBvd2Z51
jg0XERk/LCIvGYsi+F5Qp8mil07P46E/roJygoxlz9Qi+xsYWD73hQXwcgHdoxA0TsQ1dOfh7++N
MvIMRzTTa/i9/G3qA4QIGiPWyEoNJGICOSegmgUf7usORbf367RAHIPmbJdKSUscDAZ/lsgMYm66
Hf2Nul1ATVLvSRAOpT913J7PicatRXG6IYTvE8NqYc5UNtNDC0xchc/CHGOkJmZOLdrarIMmoXND
V0jQsjuq5z0nNskBM9heTi/f3+Ptcw759DJYkze5LU56ZV1e4kaY6nccEG+R/Rntpm946C8p7nyk
cml6CCsAeP/nUJTnuoFTeaocyW2pmFZLkJhvZMFvFDGkFHuZdaRToeyDcTLvFwaVEXM0xcYL6Ng0
5KjDzS0eq91qsLtSWtM53KVoOv17+muWxBKZE87xvDcEyR4iZ4bllM9Rt4wwKVJdaolHP83TlBcH
A8/c3Mymk8eNWkfXxxsE7wEgwW2jOvVPay0gO+4a844gupL0F/2RH3i5qQfYlJnmGr9VN4D2SD9+
xfIhhAeReKSbGC1stYSK8p431yi4iDegq76y+To9fXi7Nt6oL1SKCbK7mlNHd5+/ZJeKe3AV8/Rc
76UQrXuD3RLhUs8rv9fNnfHJOxHB0i24AXS45XY1nHeiE8c/oSG8jM1I8fFW5CbuuGokdHc03YCu
IwEP4/JiaxAs3zsznGsCZTSUfcw5Jw80ymAQkoqtljljSZQQ2U8E0+8xQUBYTCZYSD9jiijMLumY
WaHZ6qccfTDFj0qVBhxcQdq5ctaUTZfzf7kMMVKV0aalJUSD5d9uLp/ec3ZkKWp/VQtxCQ2BITvU
7Ao8XwTk05+9ZYPpYsZxL5ZcxD1a1dpr3ANPbcOUVVHDYIYTI+roQ3/dsvLXRX80Vi59rnCa2TPV
0bqRGzUfsyP/6ehbvrVswn72tkET/vNiQraV45Pdqc9E+MnZ+hrnxbQAloV+dy7FCnb3AmpAswFe
qGSXaJvlM1b+hxoL+l0a9PNCOWzfgSuZx2lPqcvBs5Ubzjf7rfmK3nW1/lSBUi/xUS4rOP29BNkc
VjATJVZB3UccZMzIQva0mJG3XZ4IqGe50q7wQt70uBodnZ1U4effGqLfuOD4VKYzOMMqUJpUzzVA
+MyCkz4yy4H6QSy3MbrUpAfguC9BHd2G/y0BYcuGJi7edfjPhrd2SGi4FpRHOEdzgnxeWA09tEnh
CYegWWvSiwpUq+vHHeJ1VAHcqpAQToZF7W1kBwknX0P9y7BQH9b6HnsfzYL+6MC18gVAmNvblZqB
kEj9r4Sav+1RbG0Lm9QVLBoJnQLIJ7IJthH3B2Hm1YFvoszDhB3sX7RJ0/Xa068d79MoWvimwPdo
jUKuEXedWCH5eaQpnhDjIXj4NTKNFdNhIvvEwqagxvTNtGldxF6ZgrMqO+uvTm4ndeZS+HAWJwIC
lOIkinuwT7YvtSEToEbnYHIy4kUUc+wB4JNysl8jMFq8Ve7QaoklEPZ0tahKQu5Ah43as6ESyPI0
b+aCv40/tNB/vUN//2GwANtzCmvVDsf8oc6YylvF2jmUuOUVoGyKVsg5PMCywLUccZnjOIX9LIQQ
a50SzGToD23dlVaDuBXi471b9plST5dxBRKf2XJC6v0t/mAAqg25EKt4CSRpu0xrYoaIgdM5jW4i
2dXoc1J14qjEqMM17O5nPhJwTeuGl75/68f3q1tEflYhcwMTeyXdSIvwRcKswZAyLoFLqH5L4rPU
4LYvJpXJ61s9YGKaLm/fn0e2Oe+QaXzVpT8nqAX6o0g5XA/12BLlMzt/aFiA79McKy+QwKhoFify
8WPIHg9eUr2TSXqHLQgzePzF3kP3e8m8QIOKSGnDGfbTB1P3Z+SCqh9E5dr2IcUALOn4E1rvG5rR
SWqtwEfKruUgOV+Vi313fDhyzYEpWoJdVAzZrnARbwcawARCRCbZ99iwJRWo0wrLs4UfKlNQnQoX
1NMU8FwhltBuJsfioQ2x08E37w8DAb6ze2EoYoRQpAwEgUovhMMWL5rGaK/JsMaP8jahAGUHZP0C
72vwPSx+/hKrz2peLGLcdaCNdqVWBPplQv0WZnmNZUi5ApivOToLOV2ge9orMhOeXqCHjfwxLegM
6xfAhhtIVpyNl00q4fYtx1TF/x9HYcMi+2q2wSdhgPxMCu4U1LzA7Dt8x+9dEhJoF8a7yb8MqjmI
++d0BSEzXv9RqhUnHzMOCvNA7DYVc1hVRnoLT2YAJ+JuyXE6IWq+vMmgztzTc5Gm1bfN2z3hj/WO
NvrsHPti+fAfwte/pd5V69r4q5J3nF9D9wfiTTKBSIu+1g/phSNcnsM5D2zsOWFyRsEyeq5pGw9X
NHT/z7SKlYgu3XPPGFuSf4BYZVlrZiun2ZqyS5OnU1donr1kBfhKuHssaTxioinUYCruZ5yOpwrd
HeWoPlzRpl5xbYg2IVOPt2ONV4Y+AGOwGMgqnRLprXmuLaoPXqpPQbE2Xb+UIudasIoj4r3fwcFp
e1wcxPmiLBNsH84b0BH5+cylzdx30159m7EPDH0UYB29C12hWgUmFcrzZlKQsz9XcMw2Dv+UGJJ7
nQ7RxXwH4mFlu8LHSMHfsYSDlEVw7CZWMsGM3vbWlg5oCx1ouhsVS4sEUyAWQ2tUHlqolK5pJy1F
+dTLvxWPEmoTB7iVv6TgOagbnPV8FfZnyfGWk22+1UdT/ehooYH0QF3xS58mkL9EB1oRMenMQLBr
RpbZ9zyqYj6o6jwntC49mnndCrdKwFpsNS2XlcHVT+iLG+oO6aW5LGTuSgK33uF0wXFwvaOtHO1H
4odIYkpFn1ynptFg+Z2vd0HDsJoVhtxCFt/6mKSfkJJopxw0anGrMB5gZoTVkSmJxtKcJIe60HV7
mAJ7USFO+nueEJOZetEgwbVLVLVwA3oZDeYq5XwvrWWhS/oKIxG8T/k0s635F7zT4+O+XJ5y0H+Q
2pDs/wjKSdu7uAEsogPOQvrxJNtj4aroH1rcBQduBmn3OdWCb1Ct1FdGzuGuJwIz9x/yIEdHg904
yeMzynAOtGHmG31HpURJAUoYnqM5/UK33prs7FsHBqh7uTxJT3BrODha9XikbRmUjiMIePib5bZi
QI1+kOiCTzfKeSvO0teEES+qp8zdUKd9omiYXE3ypZ0UGj6OWM0bW9bXLqXSY6gkr9TTRPOm2Fwn
KqPM6TxFtrIYDdDUj0HfcoNT0zpF1Nq93uXxkl04DmB4kHXWsjL9njh9CbMAo49qlytR5PDrwgGS
vYO/ytWJWlyen7MzRJbwBv3UZcb3Ji9IWOJe8PmipmmwcCfW4OTDWWf4AcCyGXBg1tNZL4rn8OB2
+0vPSi1mAKQ4XH2ZW7C/0EtQIS1PANV9ggEp5Do9eTSD+pyC9o2i37ePbEG7GV+GxWgX2g91Y4pv
GUfpAXjbxsTs4sC/6PxZ9a3c5QvK6CSc1I15ohIc0miLAawDregyqi1pE763g2wQqkCPSgeCugZw
FetIqHBE640/XWPmp0ItjHa1OfkZiB0KaxWiNrDBB9/EgmD2MqHNE50OPe3Jx2irKdjnfPWAxbum
nClEzA+Ntqsydx1vEmfOYPUI9fKPD5+hl/1C0j0cmecSsVV/mL/yJf9vHweuht+rxUju0bUo3Qd9
2DotD5mKAOShXe7ugTOeuDRVtTra0Qu7kF12XpYM78rZvfQrR/n3HwSpVjrKXiAOjPjmdM9QEkW0
uF03wWyD6vZaHeH6owrnEkQSIRJY7QQi9ZiktmKmbEAML6cLrayGhBibLpTJmZsoIShJjFV+Dq51
xf1F6xmQIthUuePLLTxARcrR4rEDwHRVQvhbl66hcoA1KyeIrfxKm8pR9sJzM/R/AbgO8ELUr+e2
gqDkkFn1NhI/5l9YPU+TSGve0C9IJwjXI21oluAmdEgV6fhqY3Zrubnhz2YUHlrE97vnHw87632h
iv1xoWI4lhmxi8k4H2DnAXrGGTxxIoXzHvAVvr77bXPihAaMwo4yjMw55ioqPKd5uhaLPOLmDsh6
QktkzlBjCp24Y0xo6P8ARlCwfMbOkKtswGQIsMGHPR9SVPd+bf7KmuxhbXSutoqxyiLv0PUA6Vyh
L9fAw4N8E63aNpkMBM5LoKjTUGwK9XvI6iId2Z3yK7Jjv9tZ8HRqAOHXHBomh6+GaIvrxw4yyAhw
uALmFVQETtZGxlQ7gzEXdqcL78zY45FBC8+akIc0/FCgTT1CORxdM4fjZh9tDGtKJbCu/lTM1R29
dhjDTfCNguliD4A9NL/pdRHVw3cg0c83qxIbTOUdgXEC5lMjsODJCr/oxkN5V8gme7jOX0toY1lr
WxTOSv6109ktRiygSUZzqA8Jyg33SNlISELovNd7UonpPwWZ9VH+I0B6j8ghz5XgBCcTjt7+k4tS
1Vv5Mc9N94HCI6g3fjYKiDykn24wzdfvG7fEl1PjRqeFybPRbXJ82LwIBIBWLyWZFKv/z+hsWo8Y
KXinVchqqegGT650da1d7P1C25m8GMxj9+HUnwdXRXxLInMfDZms8vh0lF12QppvmvCTmrKA29FP
8yB7GLGYvP0KI5swNP65+R04qvV0UgGjThbrl7dvFb8UygYm0FC8grsKwWHDnepr5tjfPMHfNOKl
qlu/1kDH6U63BsbMIX303nN1FLOcE48le6JU2gVVy+16/AsfXhoiRklCSwOn1ZX/c43Sn9Nt8FGG
vox2V0Cigm+GDjkecYslZr/pb1a0WTDrS7+yplYKlMR5Md2FPbUKg+gr1yMvurdLgFDGJ0b2cVWd
U61Z+GICiqQd/HtLlC0WD5iMNpJgnk6vCFWlIMgrTbhVSXXAbjuvIUFtXQZ5BMSOWDwj6vNfh5mN
6zB8a6fEZBbsvl66td6iCt9gky/wQ/UjJObpDiGFPXoQVci2RX/zACKkoxC/IPU7KltioQJvVzJu
HWJ3oOAkYR6R0LfWB9xwsnQF2x8VfVErPVTqQDGN9WEc7Jt3MAX8/sP0Y/vUvcHau5zqwr9enuzP
Su2I2mJzD7W5wvbGR4FGdiu8OuW27MFgYeO0Imzab75fOHvuLrb8YdyOZA9OdpkC6jkLkk3/nH21
uKGptGyTmj2DxJaurcBsBJe4oG3xciyrh4b2mveLwvK0y+si5MJwjE7nYDTuQl8kJpORoWSnPY1b
l6WIyzivf7X7PodnEZoPfi+DNFMm2r8MxkxtVx41lXbQAgFlwKI9/E0O9IYVR9+GLCoszEzBfTUq
CvBTUkkPotymR/nWvxcd1RAPk50ajawGKNzp2RWFrPD6DZKcapjYuEEy1geRkgX/RaZCF4bXk6mJ
zig50ktDjwb4LcjqLd+2NLuQGaCGWCRXuuuXB6hNzeeWOa65nRw9su0NvaWATC68CUAkjjQL9axz
aL65kww8bSLvW6CDpV17TJ4A07MQtXUaPCDgpLIj2rvvxx2/VMowBX0tIWMwxuuZbrT7ALL/691h
G/at1LwAMPpT9wLLNJEv5rGqC8an0W7sVhgaQ7uEPGaczrHZLYB7vMYYjvKUBKk34iIPHaO8bhL7
urBrIpD5c4RlTw6LmFkq7rmfXKz8R71/H1l4sQ0xI1FYcixAx8S15DNhNZHhUjd2g1K/8Ao7PQi9
HeAnAbOEuC4QJY7eC8tj/wal26OHQvUVggcCf1VIb0zm8hVqn4RfDrbH5uYkuj9D0YtYRdHwsEcn
AfKpxQL+46L4DskRrG0dAOh+qZxVgyWj7Shokc+n6WThupvl/X1J1ybMao9CceTIV4bGZkeBMPNO
4Y0i5cAYRUcnpkEDPL/a10V/6mNzkk/IyubbwXpP/nwFChY19Z5FCjWZ19Onux7z7IiSzVNP+24Z
e3HSx6gT3TTKl4rOxHOSlqAde9zZTbTZyNa60Luz2HH/69LToxhMurAKba0wCoahU1uEzL6j18X7
iIOshUhnQKq6HwNTPk7sq93S/nzAWZX7pt/+DIw7sptZJlwy74LXYtcsgpNATf86C3NllKjqiKaY
RciOfOgAoXYXF9QaoHooyiQPZ6LHEaDWhIDHW9TJVV2bQDqmv79iPQlWy9I9zOVwE7uqIC8ea5Yt
4ZFVS4q9Nn7VEqRg1aT0N9W7i2uzV1V8Or4V/zgNRXffGBLzMEos6Jhuv8LIDvkjszVx/hop/+ma
IYYUNAZio+jikSo9cMS7nbPl2S/77zGr0ZNolQXzrtcpV3Zf/TbnKyLzSSJ1grv29H/vIrhz6TTX
oWMQGNt2PxieM6x8qRzBlnoIWdNQouBTK2oDDLb6Llffe9GpNxc8xYDjamTvVmTZDDaRWCBHjJUj
hG6mRCX2C3898E3gXxUUDiIglVqljphQgGGt5/p5KLku57eH8MsPLLjTnYq7/Qc8n3zr6oqcWh7m
u1jiWqrlklgq2+6Zpe0HRJryTkL5BNLbXfi8+Pnei6Y7HWUE0un1WP9fjBw9L8b53nYs3RiCq/O7
JtiJbVIlrpW+SDZYy5O9EZKgMqm4IEkcC5fiMoK2ui6xZZehv2H5DppZY/nn3QZ7vszBxt4J0ABW
ULL7l7Np0dm1TxV/9R8YaW0hxnF7tb65MQilrH1fLzkJFZ3qkSlJX8/w1jWFm7sdoNP6kPX8oklk
DLARRlA1kS/wBV7wK+MEwCpWgTMx4sTk/NdlLHCgmYv2Txj4VoRNZqPqFb4Vb84xGUZaGfOX2yF3
eGvQr+C6TZRAYUM2JoXQhrxIm+rlqT27vqWdtVw7NMEwEbNznkIVm0R7icad19372u7nvEM5FbJc
1bGMxvwG428MOqK/49yx3pvRPYry2moxjGLkgUoRJfzEV2yeUOeyoKjFT2JOK352hGjPtwTNvDLa
n/2FOb7uiPS9exmgzmlkBfqRF4N7Je8hlD+K+0iQB6rexHb703n4CICJ0MsHq3eYhR0nIyng0fDJ
qcJosTsuQQSv2wj3R73M3g8ctKuFup9/c2986Fw2k4IV5MoN3Nqr32cy6b/DKKPXE11AoCwieEEg
Bc54NahtFnNhAam2NXloyfF62P50lHIz7v38deh0SkfFPxfSaaBWk/mJMcFS9xaqr8bMAc+LxmtR
3nJ0h4EoV53yB3rcIYns5prnHijReJwMQfN0FXEyrXisto+Z8l7JNipz3h+74ZhtQE1zezSL+aIA
HX6aLYttOxWZDn5ve8RQTHdFB6Wt4/jOnJq4b5l41E6SGTRCFLJeQF17Wn9xc5p27GFgmF8gfyG5
j0WRArf6RMlctm/TUs1CgQVGJiTp/LzylAGxyJz3BczBEXaSgfGkbMLfSE/vSdDuOmeQnPr9YpdX
CUM5WKoomwhAcaW0mTUwjnC37pzUIryqi6f8vpCoPjZVS0T7AM1Sqg6vJbIITafA3JSpnGnCs5s9
IlNK17YhBB7QOozp7TYNbka63BdD3R7VAVpL27Z/zHCkE6D0SG2WAQSvV9Y4exjz+bNJ6zlNntf7
ORcm3w5mzFBIwaJNB0oUGJnk72hDV2OCjKWvckLQVx7LllTbfICK5YuonKHDgXOVetoq0p1GtDoq
/WtKWJSm9ef76vYb12amYyOfjXHXJy0gV3e9KZdyLIioLUIJLEKkeONfznkhrRqvUNYqx8nhy8Kl
t9As/2zyTuDVP+wKaFqst6j9rnvEDGXN6olJuupVSBMUaXwINDoS+R0542YIKONp67HHB7uhDUIX
uJRE59J2XgCDjV3qnkIEcmd66xmNN1sXaQpTYyEEEmyzL/pPyZiBAVOde/tgU9AEFexHFpJVSVeg
T6NXuONGLKTuAdi+cN4j/LpTkUyWA5JEHrcaD/G5HOA5mKmn5E51GUtKIoygbx6wXyreY7QYGEuL
02BGBeEk+MPMVOMSVuZbizVRDGJeC0VkXlvqkWgVLsr5ZZwVSvqfNNiywiCOlpbWQEZ0iNfnHY+v
zpbF/Un9Y3nES/l5IO39rvR1Zeo6/jZtova5cd1T10taBf6KV0UJZImafaI0tDEeQFGPItX+i27+
O2fpUh0TmCIIJWMP48EhgsgCVRVZrsMWoIcvOSK3urZdjM0RtCWCvqbOVzdRtFTiMRLtIzP1WJyL
bzzjeufRPb9WJjnKbTbM3ZYVdkHaebJiomosH4sRdH73kffgjlgtrlExw4PhYG3DJJQdPbhhGChA
kqEjodvKVj8qGD/LPpuA0D4qRWtS3Zz5+QbLcxlaCcFIcnjZbDWqLFSfHe2/fQ5pFI6PuQjiOvsY
JcvZBVBUkWx6uH8NZ0VN0gXnkBL/yFs3bG2P7zO8G4BjIvebG6BMSf7Efd4fefrHgPqryv0XHo0y
1i58X/daB59F7iBL1HxYVpbAh83ZLPLriEn1/8DYIui9XOe4uVrZlkv0ra4aSyvNDTF5LKnqNGG0
9HWfnvuxTKEwKuLMA/GgPI2RS7a+fkn3JvukvQf1Me2Tr3ZcGjRP0fiJxJYLKuUtZaVhH1ecjlZU
NUzDjrW2jCo/4KtWrMBZWpc3wmfGWR17NxJyvoSY/2hnMUHybEb97vW6k/Wn7x8PM34pEK/SnRlv
RNuvFQHNy4vDajsQC0GYaLp2y1lszHYT/GRhf6/LFBis4bbsFJzEv4zVvUUCtOmbu5CDmLHumJj5
rahIaY8GpjkTfIMr2TXFdemTvH5JkuOQ+PFBfSehjlae2z7EQ8tKADTebcXeelWYpxZaPik2cgdr
ci+9BCnIRkbglkD3dsSvNXWQfuglLfWbOaKha7+hpLYJkKbU5XHz8BQqn+efgqEGYPln5tIFB62J
Eu4NjJ+aNOkRv+ncM1GrfFBoUR0vTr+Fw8TbP65GKxDQK9Qj14DnXJHJ63jISU39heQrnxi26AZj
+yc8wY5aPaq9GbUnM1IMxS1apNRtwJ/SzbVR0w4O1d6ZrNy8yVXiIUstS+XVPu7925SUkVwDD+87
b2VKWFxb0ZXQwL4debyuN9jgPnA2lKRY+BvsZJqznkKCj9CjpKkpfqz9eGYwANlIaUVaLibQq7Ql
cyDvwqqe9jXWORqpM3iD4QLU5eZGIVqnYAAtUJkJakTjyyFCXiWRtMYxYfPo38O2Lb5uL+picE+M
FmhIBgthrhr7Rym75kEXfVhfcMHBLyarFcKewxqVFz9wIYLeVk6wAvGQtZjemTi/Q2EsaDh6zCbW
v9w6AERu0d0gpNwP3+g9T1orUPT7Usb2EqGR/qERX+JPCq8wHKH2U+F+hQEdWOKNVQism2De0Fpd
VquL8k0mPqYuOCrhxU9VTSmN81KEeJkmntxM+LE7Y44kXjc+bPNKcLdi8QyNxt7OVE71RAhmUe7l
lEGr1c2c9unj16gjT9UnMohN3Pn6iTegyr90UH/5EyX4oigPuAMtcIK8sPMBtbD5PFjTPNotrZpU
5YsTBYhZgf/N69HuFOXZFj48DEPDztpVeYGbWFdmM4rJwvMwQTSW7z+YzJ1qrXjRa52FLiFAKoef
ubNpISqR/XkL/l2yaxup0qhu8w1btpHTYNVSYauLpVg9MeYpwF78GMVA/nz8RN6UOL23HgTqpQja
/PieAZ06i4A/H/Uva+emj/tsPUWe4thpNp/qTfdzCq8Q4OpFmQ2Aum1MBajPWNsE7je3MJmkofDR
RdutObANCjinkuCRVhFkB32hykEdV1fxza+c9UNPlHjjWFIWu5ihf3FDPgHfpI9kh0GWJ1US2KAU
gKPs+8GKmcI2D4cbEcz+0y3VKQpzKfrMP3u6whrnBM3ByAg55iT1kFTxzV4okEDHCv6NlTkJLx/5
waEuseMYU0++4NWgck9BqVMGeVHraUzXLCe9+pDdYQNq8/n0/NfDqMhIdYEcIZ2BPjDlFLDcjDl5
VsczX0PtYNmbWdiDCIeYt4BGGapUpMsuEGib47i2o3a4bj4MCuw31fqK3c5pZBSwYX9ae+YYnXkj
xreDE/4yXortl0ycbWtHKm9Ac55oecnKVvhDjhSQlHSPz9uu3/xXSU0xtpQd/Rp4KOXRnxBM4wCl
p4xv+ouKv/+wovRzcN0c7NE2PO93HV/d35F4l44RRubnFjG8C9uP4DEJ2Yy+0+3/zyGS9Z8KcFfB
+Mvi5U2JcNXY+lJQsQvXzGnEVysZAxX49oNgvjwpFPr5CbjXLcSF8XC+OJfTzM2HwLnu+Oy15Fq2
QVIhaJ9cx/sy6ERg9spyJC+UyGXlgnsfb8IbbVqjDAL1WJBKQ4iBnN73+uGVsm1Hkbb3Et6YcfcV
gmEEM0ejVY8UZOuGHBCH1k96WZKXrGqUM8FaRRMtWO/K3eJ4NIH69s+tHsLRUspQCdCUJ9Nc5u78
4g3jEGK/X2rycOZ8ZNx9myfNi2ZDL+nQd1tQ24HszhorXyC8lVMAKt886wqj3USM51UlrsrOGxvN
AcTJcQZ43Z7mcwVuP+QiK0RsoOE0ZUsyXZYqqCxibzTHnRvDqaBcsNkZB7Zioizun0nJhg4wCoW2
MfFrsoEgsCo4epFQWT2UUTEgJ7GT42K3K97JixA2rlUURCFAypQT505Cvfx5eZYzntXvYQ7EnVp/
qpz+QxqIr89TuIaGj6BmWzcx7nrYmpWgiCndPtl1MZtoDRjanIf9/VnWssDPFGF2PUvQ4SqSyXPW
RFS6+/OJ+PRp5VWRAVeyEIzAJjSEUkwTW8EogIfS/Zn5tfheminbcr90Wt6kqUMadpd4QWIHwuQN
Kgc1e4LLjbLXyFHMnNQIjlS17wDb1W5AryfIPRWmhGEnj+38Z2sLZfp5Q/yfz2i+UgM9Qn6dioVv
KKffoEjxqqL1DS+SO/eXTr64C2DmDECm9Rb6Ti57K1lGNC2nqA4gOdlF0WMiMVv/rzG48vJrDIWt
PjyPiiGsTKavrU2e3aDYRHuuv5UbjzVu3dUdozdt2VNbaG3NeBDGEGvGC2F5TIZR+QWRQoSSvNqW
taArLaSM+be/cFTjMJvocfI4jA1I3ykKJs3vJa+uX82+hNi6H1sbrm30ffIG2/kA72bSK6+IENCe
fSxW6l9a5K5ESLmGzqe1trwew9UP3VriBwAgkL64ou3MvvY1nzP7weYsU+u59fi5T2doz0VgZIRe
jCsYV9FJpiQKLtDB7I/mJwAPKH5BwVy6ouPyUIllyN+1qghyNgCgRi2EkJv6Rg10S8syFWgM503b
+S0xGboqdWI3zzSBnCoyFT7SZYxQyJ+Z3S+sLrxzgps2ptYODpYvH/2TeONlVvCfrj+8XpSkK+tM
c6rlFqSRDhDMlcPtpKifTCf0lWRljxYufEgCL3tNnBPJEWEn4vD7nSEJTwZoZ7vSMgkQAtdVv+cN
pYGEENFKEbZx3s0IRTTdx2YAQtRKlRSm4icud+4k0aQAR3IIHbuhyHiBkWmYORwq5tXoiJ/FhvE4
KAD5hlLx3GkiGpAt5uMkTEzkpOIYHEIL42ZtL3wJDFfXvZqq8DWH+WzN4G2idKJs129U5x0XL56B
OXb0942HpBjnjt8jbU7/lY+Q/UA0qEt1YhnlwpBD07DJ4eZy266uMnkhEE1deAs0MW6yTucTFlz0
hHr2AqgXepy8e7o9GGAUMRyWp4X7mZFXjJrWRt2URMd5O2vsABiDoTZVgrHMcMEibzaYvx8SCFYb
SJ7Rzhkmm4ijTgcctPt3c3+lIX7uOuSCtCef2PiBkG/KqnAyR/B45MS4pWsMHKS6amHdKhOkjWXS
rUZLBo/T/qSVHOc40PwExT7Rl45Ipw/3j3N3hdhwZAN3kTX9igU/LRQVgaC1wgib/cjWEK85Djx3
4jQVztewJRvqwNT7ytREpkZx419hR2p4oTb2MEvvlNbw4hYfTNTDwWqFWGR2Z271TYSvpzs47Lcy
xFcX2hB+RZSkAQJLrpmUmkouH1Yu/i47DFANV2CwFci/A2l+SRgd+NfmTWB+BSvTaOptsscSTInl
tm3LV7PGBIqhW8VQAkkuWvBaOt6kqjmU7+H3qvZKCoOh07mmpPoe9jes9k9ACjpDE3Pvnq2bnJgp
MWKY+stpf/YZOZonzgJpShuOfAh7lOiecndAZ7AgBQrkZhS+APqG+9wcbZU9MgvXEYqd6AoenIZP
0qDhZUMqYFWGI2sFiBblCm/SVTIlWGuLgmBujAogi5ke7IGdytEnwRDFvdVy8Fe4/NP0WZqMbqhc
onVCoCWi7bJOGW8H3Q75bR2rPUb1RoEMqX+cClGoYJ1dQoFwlkbY1rD9N0/NbeB6JmUXscSPlfnT
wlLwfmsIrBTdvVWNcQlah3i7kDd0T4PC8KEkftCkTNMOF8bR6zrnt5pVTFsQWYLMOY8FphkzR/WZ
Dc3q1K38BvqjObae9xVo7y8I+LoM+Tq41DaW5V3UpAoy94fjz2i3Zp0jr+djf/cmsIDHgJcfLmmc
D3+iuocDkzKVW4J/XaZTg7VbEG/OFQO4KmYsjf052bnBhWkNN/XfyyRZ0fyZ7uQd2e2Ehxb7zaIP
D3w3x4aEdIGxINQlLOGBNxnhV6QK+O86DfmNIGi6RKPmpdWR2Yqn9vMX3VDF5Ls5VmG4wNqvGPXG
OQuqbDNmSfttt3lxz7roOzqEmt6Oi25E5Pc4aFfiRQk+tYe/eufuTFB0Og1C8j/epNj5DfFkjJPi
IQREAyNViZKKlBuB5K/ofHDQg9w3WyqGUhfY3L9BYJfFuk4GnUNFyNEDHWVPae2SEO/EqA8oNVGs
CoCMiOm9rYJytD3X0FKcTmwvGQjLK57+GD9Czrk+Qi/PbqVEQW+1SPTrxE44/I4BFhij4A6U55/4
F5muGoGOn3AmLh5LhCLBbNMuzsujzh4qLfwvHv52NmTIqqjMDZlgIN+mWKaZirmh9dIV/DznuPSG
W+JpjCRZzAHP/sQrFPH/bWXuMrHpL8T3g951PHNtddtRgjiQlFYPABMkNCxwJKzMiLltMgJnn8dn
sE4wLf9kLtbHoeq1Ap169JQ7Cw9eRLmox0qknd4eIOU7nw7O6rXAIWy11ZKLQqhCyId1HnY4DpbX
D5odR7oEkwGR91c6jXzwfNzZJY3iC6ky9FY1E3MPzmQty7thOBOTz1sL/ZL7OSN8cjcPBe8m64g2
p8BzcRMbxK/fpTGHA1DG4eXcnbvu53EuQ+tmi3CiFV6m14U7A4V1CSfSUtCu5gXEMC/AL6kd+3WN
uA/BapS+XDS5MTt3ePiE7wkrFEHlVRTdW/3h7v5FyKm45tufZI5QmjF7Cj2i1BBJw58nm+NrqAYG
ZWib4HsWnElb6o4tM4q1KI+vDQ7TiqtV94WuxY3lO1aJ8yJX1iQ2toN6OyDEsSjrpggyf2ixAX/U
tdnz+7+3lmlN3DRtzZN1mC4L7YnpEjYkgvoJvawr9urJmOsYfP/LX3G1vxnTugme1B5kvJTFHRVV
oY6eoMZJrGipVr/uPY+Upn+nKcAO1gskRREWX+fsXlnxy0eqtTtDRP4WqCpQrwJZW8N9fG297n3t
lwuvA0bLh4mcrVi9KmTH81oBxzCmqW8we0noJpqRo9VMV8P3p+fbLDXd3AgKj10RkgQuQSMEr2lI
4sovpn62UpefpoFLI40LK3TGHfbMeZ5IpFEsSRiM9tK06sTEpa7U3NSSMwT+5lG0JjxONV6+4Ua8
ZtLuc0ETmsAlRfh1GTc2qVDCY9nbGHZnvhSAIBpg/c2TsZ5ZEWsLbGxpg8YkwlFskGNdbj5ok8sP
yXcotj5k7aeircs3pS9XqAx2X9JuWoVvX0F3skgR+6+UIIY1HrXhrUOqfLKnQbq3m6nSlbkbNZc8
Z/v0r4AVYxXO/VPs35tXInutI7ZzIrGEMuaCJMEbJMIp5p72Hj3+nqF/RD8mQXYDV2Zg+hzUMDQX
kOpzE0TRhObI44gOuGklyl1juwyHcapmmYcm/OYZYeSWPW8fQQ+Oh/5yyb8MK52E64SfqDQcVU/k
8nlOntxdWoyYspdXId6M+2QTNuNQ7La0aIBFykzHhg/Aet7inYzDtYbSFoK+KAgRs76UpUGaFhTn
QQIIuA4nTTJpuRrfxHH2WNvx4Aa5hPoaJRt7QVEFSgwWWSEj+ZHzAbQ8zJr1uZdIawv7xia4Yr+s
zzgj0Oc4Rh1JCObGfRSlXERbZzKZ8MzXS2AP1jnYU3Pisqm6DvKyWOu8ojnpDzOGEhl7i1a39n8A
qAUeqWV/M4+xPNHqET+8EqBJ1cjUFusPhYmgmczH5ETx4GGwVrnk6ynr/RcvRzK0ymUbYZ+xpqRO
y3GvXhANwbyzAN9NyPgrTksiYJ89ZOnE0DW6kab+gdcTN8uZwlJjWDTAAsDwrlLxL9wgzxmmgml7
xC+GWmx4EvhlytHWqWsPREEMCqSPMPKzLfHGq/VZNNgdyPgCck6DxuHRXYg3i+kvb1/IDaSmsnZm
2oz1OAt+eWUNsDcxfJndKSW1+NIAf7Wg6h2hkJ29OMpY3L8Ic65oCgpugREVOi10bmDzWmJ5y0+R
fwE3xLb15o4CKBvl3/wJ2Wf9ERZBFoVqX/EsezUDbgD+XQ9qEiioUa6p8oRrSLqELMhB7M6pXAx3
8Vx7Kle9btYcttVz1uA6SS3TQpXmfI3iiu5qWo2h/aRXXM3Pn1jUMw7K9XdVzb7G/ZSUD70u0uxM
YWP3xdlN1OsX/pG3xOLpjPicws4mH9kkpU9lRkaoRGpWhs1jEm8OuHhDsDVRz+omappMBAW+IBLx
5xRiamT/iyQTt+9K1j3yIm1/lK0QybHZGI96QQSbIh/QyFkt018CiByUd6EwkKqVyjmJiz3tAV5M
g6zj0FSHoHxyW+hvrs7WPnLt/504DIe8ffBlV/Vrg1+831QQrY6Zj6LafVuvhLmpOwNfV2F8eGrR
PIwIUjWVrIC0+VlH9YhBBWrO04ijIcZNfH8tkRoFtmhdAvI+0oZ13nyAsDAUoisnxDFl7s4OS0Rx
HkalSjGtiumNyjR48Il0DNAO+MKmldnT3mwaL//4Sf7BsGERcUWtEciMJSR3KfKulBAV++PmN7FU
/8S/IgYY6fMihML/+xQtustR2y3wwc/Zy/+tw+ikfktzRunY0pt/1xW/0sEpWDEn1g0KTANNBsSP
oNZci5TaWg8Z9GmEazqJ9+b0X6Uggw/uFudSHxIbUqNRWilQGEeKMoagRJQgOR72RVkEskrmQZmk
uL9ryIBWMzL07r7t3crYy9tbVJiRIXcuYrKdyBTnzoFO9ooDqngaE0kaMFy78TrbYqddg0rm0cxl
FhJlHQ05W1ISgxSJJ1eIp5MgDBtLj5rj0fuwPG4+aQRREJRVjvnz+An4qi+ReADI/0opLMu68mJ6
ofGB8/yGN/OszwY3f3zUd99+fT073M7kfKzY6pq/JneE9bomYZJE1PzEEt3lstNL7vrNg05/H0Ko
AKTILn6/qf/nHZh835Q1PBu9z7w6n1rfYNiiADbbq/dko4kz/YdF5dEo9nEBmmstRSoobBYyr5ov
XPxa4Uj7/Eefy3h2dP6/53m+G00J9q5Yxyn0lxLg+Ua1t1oBh7EJPZI/oi+1cNzMMRNb1bTzrAEr
zQ1QzV3wiSlUfTPSLgobQkMnoRy16e2GnfjrKERu9LEKeFp40+BrjP9uNjsIhBWNVtSN3vq3nE+i
zE1tCV07kuN1Y0dYDO5fEJAkV7KRsLxpRbMiXHZVffbVPgC107bzBKRtvAjZBb6Ixk8wXBbOCN4I
ZmUa4EuhpN7urTt20PO3Wd6TqTgVsmfc6O1/f3mxJfNtmS+NmRxAsGh0CdXBZ6+KOr+Qg/LltUYc
bVMoRDSqk9GuGUiDU8is7addJqKxtrzvMnOrjL1N7O38MbfbMaL1GjpzxQLJfmbnoNb2ZimLdAVG
EJhqvAdML5yWdI6UC8ZGrjGSLcNp5w5cXGg//K0zeKN1UuSNWPnJeb9r1UFaiW4dyhKDMss9iSWx
Pox1T8CMj0lG1+fxMAybyh0KUcfwoEVisSVqdRD5iXj7PprzFXzgXgN41x6iaySSmInVgxDbTX9w
F7Uc8Crbdy5iLFRwGhZyBB8m2LNGUsTvtXJhq5vWoXl4E8TQ69jJI+grY0wtSxU0nG6RCo1AMoy0
C9l8EBe2aZxEXsgZFtlihGJ1pkmfJfhviR9w82z3DLZcGRapp7m+rUiY6le3ltAbIlTB7Dk/kb2Q
4nmNWzUyqohMaPdZtZvC9rgSsngiG4Dehsdo88q4u5LIuux3fnMor8R1kkhFmH0PZ00h+Gj3N+9P
JRH3tTTI9f73gK0Q2OHOXGxkwOg6oJqoWMisgmYYieM5S1DJn0fNj9VD7EViLxv3iAOo3ArZKjeT
xfHq7iM4pMTVchMuF/sW/yhC3WSs1DlxM0oPcZTceRoqDHcGBZR46hhe6a+zIuJF/pDIBI4GMVJT
uaeVPxZIud+QdH/KpqC7ePo47YNIusswtDqSyFRopkaHHijm/GbfFEZ98kiDKpyMI0OBenfWAX4f
hT+0drdtqBbipZQ2cei+kAOWEmqQZFrNsT7pezUol7sot8HTP2LEeiyZLCXoXS1gx4qcAzjaCur0
k+4RS1seJKKyOWzRf1Cg+5wkFexHPU89TVSj6GS9w21fouXZLKJ4wY5TWM8uyAD/2ZwU6ztHiJIu
wwtykxO94qeKJIsJZmBlBRc6ronu+HzxrOTOiZdy+2bGQDdDDwjBvZBZWAKpN/qnzwwnuMX5e/zk
R2DOumgHauuUvfY47YU9PWCo1BCg/mJk1JOjGZ3bnPVUXb4s1LbzQ6mYUIFuZtVIX/8d4f0H8P5t
D2S1fYTm/ZJ+7zjMVbbSG8rZ2ya80nojKTIEVS2T2M1xT+GVcy6IQAkqbZ127lpHw9hUuyI6Pb6A
BcPhmZPt13SGG3jhnFlGnHxVjXpuUwXR2UMhH6nLDxuidJUMpLp7qngVRtccx/624u+URYwwBYIp
8YWbCmm9JPVo1afmXkPipWLW2bXdr/g/tACHrdtJ93DLe5YtddzpS8KfkS215aF1RZBO4vY1fUU4
9At3WIs6tuXeb+eEahzELz3zH9BFDnWAeLqUiZighYA/sO88kfBCSxPg8YsDfSqdkdBWK/DE3lJK
l4WW+BS0s01ky1QcD8M5DAKpMf615SUCnxwpqFnM0VNAb5aOVuoH6VUzOA7E5x/VAaN9NH1oHEnw
ak78WGwmryKJVuvOH2GxkSGjE1OuUTvI4QuElym9dhVLfLsadCa8c7DdRqpMhw3VlboEC084eHDC
b0H/RBwkqNia9BRWyaQi1tvp/0uAJoUxtYw4N1OwfHIwOc8A5vDf5qwEIPZ8Pdltp+gZJmJF4gJ0
ZWDf6L5rCROgVs15jidXIKgWpmULINDMRTguVltYDsT8cYzNTrJQXKAp2plPT9rzK4R/u0ldkOQH
ZnVjaE0Li0q4YmarIP0fC3vsGJHMqKi7l3uIEbSquBdesedFiK2jiyKlV0ifmcds9HQdg1Q46F68
s8YVtNCI5+E6xV9J0zKM+1QtQ2dkRJc1m9XxUHiWoYCzsnBq1iuUHm/aquxxauhaNWS5dxvYA6CS
ZQDtmN1zb7SV0Ewphhfwzoyy8ODfiqtsXQc0qrKE1EkIDUSc04hitISLxZVV9TX7C8NR3RD7gpV3
xamKyPKlwdt9xKFgpzv29YTX1w8rARdMRAvCCFNJ5J+zmcianAMtxp83vgPhMSlGrog7lMlDhSBQ
BKo05OapR8QMNhW/JjChPRJiZtdVkikBanrywH4+Ckul25w5wKQHlmYF5uxe/x1MPkVGE1EXdEDq
04fhqZMeMGjJ6yf6BYKYn+PekIjYFiewc4+K/EyhUQTfhf3D26QFy+f4oIL2f9U/W6ZmreOSO1W0
azHf7emHX9dbuLkxqojqdhmthJf/y1dwvufVvQA7iAGURH5ZurAAeqY07XKFeWKQ6Y3RK/VgWZB/
uxHvN0DNWF7UH7DjtppWQUbrFB17f245+jHpM6wfvq1dv52YT+MMWbJeJAMenHN0Paey8P1oWHqF
Zih4fkzckZana1ETj4siBJ+4G8tgbKJL49wHu1/ip72kOv3oei/uUG9BLJUQHv3Db9nbG2VDCoA2
n/lo+kHaGi8LwB6ObFq813smyENJd8aN6EDWRo/t8iZkUf4fAXrXmWf2gkfWViyd5dQZifxelULO
LtqsixTI8QgKpwIHuDNRGb2zyL97Eb4X+of/47VXktB2vq8me1g1kwozCH5rxIfCAjKCWKvDJ009
HVUhWc6Nl88wzd8AKUwmCk/So8Y688E2muij1ASSUmqstxno3MZWnHd7ZLdBat26b+Ce2akgpy6O
+8+LrXPBaxHVkkR74fNz1Ug5Eox6880uXeqLFP3qYZsg54W7ab21+E0phPo77Lk7/oliyxAEhRsn
3dhQNz3rqcJmJba5fOZykH4coBMQ+R0508aPg450k9IJcxrSCHsWPbAg0fSNwFhog+6rmb+5c9k3
lA27EqcjWrvIl8e+f3RnJD4GFfCAlrWpiLJGjo/eyReUhnsEfqnAfYSpAzIaNemwdYpoDeLe8+h4
nofshQd7Vcwg00GpAdI8CWcA6Qyqb9wxQ9risqr7kbWiVHQ+lKtrEnANHWApd5CVASGT5OR4K2W/
9r7ZWknQeRaFzG5HXhawILI9nlx9V+WnRri8CgGVrEQS0Q32RTpTV4Fl4WVtfP80HmwR1WNIff15
5bBnudNw3hX7rNQV/7f3mqayttWD5KLS2Jy35YXVFFIRlNReyQgt1KM0Vb0iwUZnC9PMReT+68oo
ba7nVCichuWs9jHsVXtOdEoVDMVsfUlroi6USqoXQuz5udOmzNrq3DDz/nKMLeSIGd54jpel+TJY
fHV//n4yMVKy89bjFN15ww4/Tv9Wcgt267jcIA3rb9ON/CIglnCyvcojo2T++EylvSrsYynzwcFk
Ki76+ry7MXot7H2tG9F0akb0dnB8OVlJ5e3HlQ6ed95S4ciGCvScMISWNAH2bCJIVZbnMKkMzruL
SwxwWQXAeo6jnd2Ji4gudsJdkh4qzJs6KxzU2VtO5lNLhBhiHE3bBZKzGv/qq6YUqlwGUV23wZ5R
xPmirZbwszU0xg7KZPxQRDGcI5B7mGB/ntQ5DAMFHaNP0oJUR4FvO5vlB2WCCO+LuEGNp5s8b8sA
UU2tnHbLcvUAoD8+Tm1NyChOEUil6VVwKYm2ynJuFxudQqs2wUQsky8DUAf1x6W/6AcGKqfmUaa/
OiJRIuBQgv/Jjts5SZqtxXZaCc/O03wcKN+wRuqH46NZ4bt+mFFM2897Pf/rLIrpqhV8aGL2KfeW
198Jda8IhI74JYvkIAW5KEioBjU6OkWB38OZI3h6iVrM4Pzd1DqIUUXWPec5MhTDSJYpiu2cLZUr
929e4bh6qmIMFLIX2JRuyhV8h2QHXKuhnpeTURWQtnOkGPJQsmfJKHOzunhXPDhL2AAVJgZ9XgmY
287lUuUjUW4e6Ubo47wDalt3WMYZYZm7WUUHfn3J9PnjTcF9Ctt03UYyiU4DUEKmT33W6/LMWq1o
a9yt7cQ3Uvmycy9cAAq0qDBu/aYjMnpMQ2Tl3N2wMrnTXKrANH7zYTBAlZ/cCQM6KiVda8cbgD1m
eBgqa737iN2C7N3fcmwjAoxMKzdhqtBWpzumyMVnySapyYvxbiJCCyGXRdbpoE7AjKYvBk3ezZyD
QE7MFVnoZBNVRw/6y0bVMbrGBLKXVK4Dtx7F8VgvAughmRYkHHfDAZ00VbPPDWUsVhzn01YbHdpC
gpgcFVfVOttTW464MrwpaOl29Czbj4U6Gqz6rAMbvSwOosToU0yAIAF39OPtzNoEXn4b4p6BL2Ur
3F4IWcFMX4T4JfOGxq/+ZtW6++/ftahgAJ3+6uhBtsW7CIB3bGg9vYc+hhpMDDh85WYm1p+FxFPI
Osiq7Cczfkz2Ek3IqrgX2C5bLKQEqnQBSCbAQX2cSpZCX5VoY0uIfTl/zR8/UN9gBJPLvElTphya
GTi0CTm8GNBnUQOazYUb7EewDAMLEObspE6N8yyGiLwjnelM4t54UwDew+YrzAf0V5XPKEYidSv0
n7QGVmk4ahN1LoOGgGQruzcTxoradPSUyvzenfMvcR6NzVK0B1U/pL072hBDVXDKq3ZFSCYw6TGd
YhQFZWooPQSTnDMbJYzKCsB+zUxeG914zyJEE42Qj1CniEFtFPQntezP6UlmZLmoXMqPKPeJYoVD
LmPdm18tXv+s13OKYpbzIU0Bdg2M+q1Bz9zo+Mh3aSEsZI4WQbw+BhKg1cfQcv/1bpXfy6p+vMOn
trIy+Rj/eEuTcArVIgpJu+2Tgo5cFQ3muq/0NWtP1KQj4AspVwBJk/PwVJdbcU3P+oWy4T+fToTV
Tq8la6HdN1tdf7pr71PnLJzeiwkxX9XNmDa6GTUAgVWZda8ygPexttFtCMIWGRxp6OYggLT4a6iD
yA6dCZ2Pw6ghkzUYG6F+fAN4WhFrX1aswADuo1YwPUQFwiMAXaFL/O1+Z1N73BtdGODUda02QMlH
wb9VdjXQw9uRXSvl6spJniIzN+DKF1B7cxIzfD5aDvcJl0wXf1zYiBcO2ZFWQRoTsFcSMyiuku2Q
avt6iHtX2b6wl5bAo6Yl/j4sgst6M87dnIwp2ek2Gxe/4NSKRvfprhqpOnvPdHzulAkdkyYaj3UM
yqx/Z067eR4eyns0jdCbevcOikiy5brN/iezYmhOVBz+/Vao31wdKamxwjLPZUDvUrWoxX5kKZ+j
RkyYeOaD/UGw6IJ3M8lQN+Obve/EHGV9aX1s5YoIC997Y6MLp65aCNzLw6tMXrIHlJq/wFw9fzRZ
+1o5yk6iZ2IqBGJujdWxwaPtwVGw3PWMEoJZacarntGb0wD9f6+LNxdb8KjqmIWztTBZReLnLYFW
alGBQahGW7zpZ2d61r9U8AaiKaRY4v86lkTI159OFkzXIA59JmZZgrE1rXqrUay4X23Dh3avgfKd
UHlKv8khmhGnq0PeBECcYAN9ZbdZQ6DJ/W8t5GjtyvraK+bnCN1Vldu0xxIal+mErYLns0pu7XAP
8fBHfo4GpR/8bqIUpdHuOEX7CXgYX7fiy1geKX4xqB4hvUe5b3bMR61TcK8uRvy4FUOpDdN+5U19
Lk3zYZfLEBoZZle1bJDhEWq2QGX2m4MMIPVTOwC0jYayZ/tNbDwJUfk/0D56U99L2ngaqyPnSBdn
3aI414tlHIIC6AefY1R0rAG83dTImxwU41eRlRV/MRjIIJWCjhhgB16gwBNk+n4N1idiYDRnxVub
yiZFbGaauwKK7OREfwAEbOQtvobaV9JWdyxKDy5vkjuiJhBCNBjvz8pr2sae60yhM6JEjJFp5X6r
T7c6ZslMp0uLs184315EMDuAVS3DjGzJQcmYnisVMrlcNNWu9Xtq9CtySz9fEz/WUVo1+uuoFGFt
c9MblL5KjkTtwmlPxTuX4dopoeGTZ8iwJueZepFF3W38MY1CBqgCJV5KKHaceU3hjOOwEQTwZkdt
B9pTgBT0X577L/Gdmi4lX2I6jRbXOQNkq8ug7aTtpLVzhTYyjdqwYQ1paqnRkfL3J6tPV6yBli9/
ZJJttQV1dzyGAL63926FFhfAy4+Zd2CPqvyuqy7hymgP8vvLq60QANwTTiKvaD3mZ+bEO1oHUiC3
kvUEIkHOrmRUZ+UFuL2CMWCAwuc0dMP6/zFX3ciJZw1QTXNQETKMvKLasi2IL15mC/8YyNuE5wsO
h0HdiSxGdxqFsxEgz2hEx4B+15tuZcjOM2NaNhaTPFDPD2ICh/RA7RTc74KNXzic8SgkcjQHOJnm
3+Swakd3w7CRCbrBb7Ss/rM4BleB8Li2Eyr3W3r83cMRJkc/QnRV8FXj6z5THw1THdj70kVJ2fAW
3zl2arwoVz8WWGn4GkiBWaVmfRCusL3iqn1/7mYIDuZnHhV2c++ww0xLWyulj+nhSulWsaPeSrt0
NSW+FMYIYpqGBIMr6ikHkuglz6dWLyNx6DIA4CcqPlTf9USmDqFjfcxABn7RbzDcSwt+84F2yeLu
rF8etOkmxRvvp6L4gtqfypzcVF+bmJRFllwkwr0q3MCRe6SycsbGDdVdiWB17vJPG194FV1wO2VD
kmsQzAXeBhJMuLDAu+iFUUYveoZLWo92t1xK1Ni4Yejk0f08N9YjD2cpjmgMiWBjSo2z63zNQnNN
0ttQj4JgxUIaLzh8e/+5sb2dVtPhRflgh/uOnw+RQETbpLxcbIV0ogze6QUb4HwMFv8p7LzPohaf
W7st1OWok9s7W0wz9Fli5ZepdPKYxczXkBPUFXvPUBb7RzW1Yrf+R07zjZaWpt9bxpNcxTf3TDlr
wyfOsmU8X3kMbLSbL9lJu0Tau4OqMCiA8qmFxFBrh9qDIkLv+zzfNxPeQHLQnRhcwMf25KViO/XM
7rit0/9mRfnxOJ6OKzGW3rk0Fej3O7pdiNNffEq9z8WDX9VCe93LAROI09qMTcTESubk8RsuDaHI
Ify8Uhh05dz/E6CXHBgLv/wKP7yEZhcw4IzelbwyyxfeLpMfsByGko6uW/86d3wS1yHcCK5QX2Sl
9tAO/lA6xx3tlpNN6U3crMffwxeZB+tf8GP5jaa6sCz7pf64d/SgSCA3FwbCvGdQjfHTEyVIkkUM
XecuDkEAjdFIXAhnHUfF8j4R3eQmmCAlwfe1aUl3GxkqXmCmdesB9o4Fqvnck166UsprzQ1Lg1Kq
6phGIuOnVwhEj5P9nuV1W9YRPh/EUPaNWlr6R5sXLWy5BpKq2QgKhpU/K1PNe8mQTNmFOHn4SNSE
M6y9CuBRNV0lRaX4UglkR4A2qTM20gou3nsH2m2JsfRoSEXhGs/uxiFqVFYl/HHpH7ysYQdEcCiT
F4C84ZqUnwEwfOWwCLdem0fGMl5kGTvoBGbGVyS9h/CnLmZS7HCDdJQYLtY682DFJaUu9BPPl0rD
HIq8BhcPf7//YpgrJJ0NrKDKvWL67mSIChwFioZj7fZQPWo/FgDHWpk9/8+OuQCJfJzZuyAg6BKL
BtZ8PZg/gX5xhTBC1aiuAcd2oXu68RYZq4CrQlZYaahMXuWGF7TBcf9Ou+P6tR32R6qbu4iU4X1F
UJ8bsx3NjigYewjeFz2LI8e8zIdlDeo/++W1+lckc9RCvJt1gC5NfZ/bcpArCRCGxN9Of+6XL8z/
6fK9X4FibFN6nMIDozhnLbsAgmAdTjSiq/XmCXn7KJ+H3sOG3pil3vLq/UZwYYqyuiM5+6sIu4A4
tmmACCJVFUm1CRmoE6XtKhmt3VYLv0tOnzsMiJ/vZb1VcoG+08gHzq0ur98Rrgtte7f5TuQC3ZhZ
Sdej9Pttk0QYu78EiIBnyHzwLfehzN4eP6WSpftAq7P6haUij3TnxvEPD/5MqHVc5NhNGd4mGTRq
7Wz7DoTkIDnSHrbmSeLCLR5n4tn+ccawXEzar+BVwam7PU75AjghrgTmafSxN2MAsm2fWmewBLbp
1pBB40Llg9pgOPmGY1vfTSqY1cT5YvTJC7FBMt47/A1S3uhE3f3RgXjg9MEfw8TtC8LI+BkhMHd1
iqmO3BLH429AX7CSEWHACtfdVSwiUYUrwcpoX1jyoIEXjLtONzKqitEXQfELzSIcY4My/tbvmIpC
o26JGGyphY5XLy6ohUrXbjiekzGJ9sdcAh8tsGH2pvbir5Pl3xmHDEF/qgM8EAsa3jYVXhEh8sPu
rOSCYIiFidYtO/jXXP++R7tvu6p0Vhl6odhGzHpxVwSJXwihr7SV51rWRna+L1D+zx2sr07LSsyE
NDiprnqmNjcYob4TkYx9ux7aYw27jsaCvPp43g6RP68vvLc5hGoX34o6HgbYNdIy7yjpHDUiuBuo
P6oosuciQCzYaXPgxKeaFXljWM8yEewdf7jMI1Z/r51A7eUerlDXsyKOB2mwMy3zynOvu3LKiPNQ
wFtgq+s5eqn6uHGK1SHPyLV9ECRZwBhiZiHxNNTa+4/LavqhRc4JU6kFFwlPmDPCsa1qE6NXK6JK
z2oGpzA+Hl8WWRn67eVUC/tKRNXr5Gti/Ar+XLT9wzrgESG4PiDB13EAXYFWlhNjQkrOnSV4TduS
oSNhMcm4CyPkoK7BJbMOIytrDGoC14jYegmp9XjDIa3AXDHsG2liWxl/YVI82ZGZyYQ96ZtlbDwh
gIDsl7ARz/lrIR/eLRgJ14o5Z3pVIeMAj4seDhgUPDrtvKzamOB6mpUhXKb6DhtKz79H7HTGwNif
PiNYHbbvBVmMHrxt5RAIUNEdYFaNK9fCgCFFp2E6IK0lYKjni0BW7Q5dwwAdLHB9MpD0bcGWv2gH
a2DI9NMJlERc08cA+msHdth8Xyhk4FB7MV8lt7mE1ehWYvoI3jcJCjHwNidPx7FqlafdZwQGpAoC
fzsBxGp+E+fDeT6vuQmpBS9WKB/mwSyqH6aTVyY9YnCegLCer2PX67xfolaAEiCX+ui5VaNtY3V4
hoElRnysVCIx/1KEWs+PCV9FZlSKK4ByILrlbjptzrgq2YP//sh3Ad8Ku2lu5ErFwP2eTbmPycyQ
Dd5anypdgl/QPUpim/ZOLfcm9bm9HIJTEil4T07lkAL1B1C3HkBLlz/ePEZ9dN7kRlFEmHBhCn2t
IyR6Irk0LMR9aLF7wUcQmo/PiZREuP2tRKlxZDZfW9AcP0X3RbUkIIivNXMcmrTD8VTC409r8wAe
+hNUAebIAdOBBsgNc3NIpM2pufuWK7wTDgv2crQPnhg2SZYlVVUHcuIcpM9340qK9iehufhyjeJl
JkUa35Ds+15+CNRTDqCN6wTI7NJ2Xj7NWkKLopS0wHniiAPJRRCnIFtmAcQxQCaOSJK8p9/tBnj7
XL4KxXQk514I5H/GNAwiqz9MqfYFSofNrsdajXKrqmLg3IkzXLV/yHPSd5JK/OdSxUFn/BLfT1Zm
WBrq7rvPL9p5c4nx3/xQTx6pCTXUAeaW0JkkGl4UdAT3dyvuFaB6z3e2HuJS1TiHIsKNZmFaC/pf
9ms9/3gSptzIez0Gzftwkz6u6ZaRaBRMwzT2Tnb6s1q7W+xfZtBsmQsFRSikZ6GI/KgM3upfbNhi
HJyLgRleJo7f8MjA/Y9DuZNTgtTv87jgE+08MvHho0sPS1q1iFbKW0a7WM+Vtu7JCn7BvwtrFIO8
Zz2iuAogQ0bZ85ZEnVOVo0P39HDc9V8KJGS69fb3R0n+Skte4PHk0jLk2UsbyoEfLID97QH5FeNx
+5ksUjRo3sTtOgJj3hALq74USdcQYJZP+T4w1ES51pq92uW6XbXb0GUeNU8n+F22///dxWso4BrP
9BuX731U5LSadoXBWUVH4sY/wmELKakPYk1fTAoJXbDHHMXNqdz8dN5kQ+Yl7OdhH67XvdqzNYJB
YJ9fqffjXYAg/KCvWoz+jdKZ1eU8FMaIio+2ap0zNkkQI4GeuXQ6c1XIns4Po5Kbub6/YUxu2tV/
xX0s9KNXx/aqocRqzQ4HKOKXKn2YWPhY9KiwMGxFO8uh/G6/oD3iOQ0GrNIiw+qEm+w2UsGtwFI3
ql7YBsNQ6wEZyMs6rplkFCIXzTFuVu2NqcNvbAZlOnmAQlmhcf64PbDDVhbrzW9hn+iI7i39ipGP
j8WCY/s3E/dXxGu2HzSV73W9p7MlHNz/78bt6yz/Jv/ACYFyxGRbAze9HIarz/GtqKHIu2kUHehR
fSdNXKXW7h9VCIp3tOuLrRNBjKJ0eNZa/PH8BADakggHc5ilHSN86MIsk9T/mOSlRhpLKb4fo5Ll
9qjGcpu61WLCahCY1zU83BqYieXMnswFImDxR0auL1g7uANn4cCqlwrZ5FvHHbcKQ2WjME9O+pGG
8/ApcXosHghPSm/RYUrvPp7xB0/XrjM3Ad8IvPCcsRY/vd2rYPn6/yMReQT26VB5En+4yYHLuEmt
UNNoelGgtbN+hsSYlSdoYV6ZR9X11aoWwIA2zdst//HsmXIfn3E3LgW6HHfFbnvhR2AONvWzilmA
xby8rkWwsL8nTbfv3rp/Mj1ama1VHGUbhQHzL9sMdWx+DQ0E+hsZb+SENuIdbOV8R3QZvrEfIVFV
hNOSHBdpsh0pte+7vUQbmyDSuxHBsyRzVYDsGpPAoAeapFoY5bBNUsBMB6tdZFgBkkZX2j+g8GVJ
Ce5j0Tf/gYYFVk+57dujKmciLei4YY+7INqSpIwfKCUoRaawJk9vwNLVzHBP0NaQnzvyXULB702m
568ERN4Lc+kJJ5Y4Fs2pJrkW5tePK9JdSPDOOs0xpBBBBIPDi0KsSQhGldenIONqjCVGKhLKHryW
GgKXtgSe2w1rP6Cj5Gt6GvuJhf+Qkc8o8M3JiHWhGukC2UlTH6Sw9KCgRVSycJpxOf/c2fza+UXJ
ZAb0gcw26cpJteuSMpLIVnAYm/jU+OhoqD1EG+1xzrnQNooj8ctprR1KdbrqSUQORD7jWAmlE902
6WM3jpBvg+WHSlA19LExtm1YXC1ajA2jJfuzaaHZZox4Qg1V7e7FY+bLl2ECBtS8jM07m3XcMPQh
6VNT9l6GADaUn3k81xMhyyaj0BDB6QL7tynpEboc9AA5apDu6qxuOT8TX3OuyrGu/UV0EmKh7wCk
f81luDODXDENVHpp2w52mpCisaIwrudTWWfKrQmvIBfF+rs/s7WpOLEkGs4e6JBzaKfmDyHN1WqM
bB7OcVe8TTkj3XusBt7yg+Fk9pUSNRRIqFn5bvHMk1GVNNTkkE1uJWkcM6jSRjBGvbb+Fmf1rv0Q
Sz2StYFh2WNsAsi1ei72A7Saz8byuyPxjObm5Vf/dWHG1GBI1thWxF2OFw34ywlyQUu9AR5GYTRn
lg64rHj3s+DcHewt9pYZ//uOsuxRfmYryo5+cVxBVqCFR8kAytdWZHhQQC2cmk0udosZfRkaEacC
RUF+zbu4VIVd3ffF2eRTY6q+COEAA1vwL0ojRaDvCf5XtAMDkysxAqmapDUVxAlrIS9MqOmn8W2t
QAMXVW9+ECHVaXQ2CqXe0tI8c2/9RpD5mkPBAbjXwbEaOsRizGnvONp65dXo98Gt7MD4ZsW8Wr2R
Lrb1dshpBDBFHscmg6Cf1UKD0tsNtcOs/9X7hS+dAoO3a6c3Gwpf7z5IfMhbs4sTBpT2/P5APFqF
avh3TtZEfvu61yQfKtXz35pPjP5xgfUNfhqgCnFUDmzgNi9l6r9Z7tc+jpBByi9t0oxSULFVkZEN
ix0TpiwPn2T9Z/KRUf1qQoejIW2HRhVx2wxUCSHiaN3IuPZbZo2TQ7EkvFv45VeXS2ZuPie9gqzA
kEEls2B2CZbJl8BfSa/uLi+3eY8DoE7GJwQlxpAxy7POmSl2rczvLJwQBwnZZ5AUcYZz8+hvns6c
8a1rWr0++PTc5EKqg+PjylArlMLp6xBHog5Hvdz2GN+2KfbgE2+fvkCsZp0aPMyEB9CsoPXyK3O7
5cSXGNJo77VOG71WHbBrTpndF8knbXh9GV9mXhasBd3ocj/2O7OsF26D966nDbpTiOwCG6bfw9Db
qUZOhHdtQmZkroySjldUYHaLWyUPWuy4WaaFU9MXNPfx8DgOsj5TM4HBjDyF7aYI6WCPKfhIf2bY
GeUiS1QIEiJ7y1Iz8Qxubf3uCHOG8eE/4jJzD57S7u2r9Gs5itYA7qvktd56wePQd+Pwubg2PlcG
3SGzH1HXcMbI4eYsvMZO2jVNFdKoSHpQMchLuKPPVsMXynQsPkAhKS2acYZja7imoc18ooroTNyb
4+BPefkFtm/yz5J/XRkIKPMFnvi/29s8U29H9VUQrYWKfsmLKCkqjnt72FWsEwNEB3+/H7AKAmy0
GoTEdWgzNxOKO9+q4jFS0qr30ygt+VHf+4JnbULxQrPlDGZ8Q9OCPp25zCmFjcvXXGHgp0Itbyfl
7cfJ922T6sgyyq0D3xxHCx/mRw/tiiNB5Tc3pyN4t1ACQPUHjexSsWFGAOpPjzGPSp3+WUQ+DRgj
6jxuUDl/V74fQAIkvn2+Jz7PCu4mvRpMKqES4PVZs9NlOGJgfeeSn5y6UfiS854jozaS6Xh3ZiRz
k3PMjqqY6OZjBXbERiVDITFd3l70OyAZseoHcCGaSUp4Jk+Fp6G+MWpWAYXuhXwg2Vh+77/g/447
9YH1YLs5a2j82xPv7OBbPvF01CpH+dJ8f8VK+xgQiP0BzufYXrcgptX/irWGVa08xFyuS7w1ivXe
D/hfxXJmefCAuIzQ6leCMWejScCU3EiQgKmTOsDjYi2FrIvPccWgyLFRBCID8oiYhJaIuUu0efHB
3kM6ZHl9OrovuKWQNHweXFvrTs1+L+439FJTjwBV4UlNdVuRfwEz3gN80ye4KxMUOVO40VFs0ff1
x2sU8HxYaCqQQ+cdtAHIW2sXCtnz1vRHP/3vX9LPYCZ9b0PPdpSKZsH+jwgArqPwKxC1/HTmQhjN
/5wFen9q4T3p59h8cecUdaKZrTdiEY5xDkE7uVqcUyNZYx8MLfIgR3ilrLl+wCzA1hVPh9bIZkhj
O1VVcm+8la5EfMF+YnzYTW6e8LNyx4/n3ACmcIKoSq1TekzeRJJyrRfg63fqjz3T/kDCaq7RtkjK
tHr22SV08iB/F9EhiFJhtII6rMq3bBWRRa+2cPJ3Yk+QVQ2gxcfdD4H3dBJsxIg4vCWNXxwaEW4c
8kwrvi3cPLN+t0MzPrzJWwv8UY2Z840zEailusfAA04ql+UUJ6ElU+y6JvbRbSw8W3LtSdE3Q3SZ
BZQ7YXkoq+ccM88RXR70+D/1QOKB7ll0pxuyL7+d0RJHnMhoJ81VOc7+jbQnQbVm8yV8VvAIA9Z+
bDwARKeQHmKi20XOGN4ifGISDAtru8TgWk+7KwdKd2x967rF3jUaOiBi4nobEHVfBCPtNHTNYZEA
8Vzpfu2DiA3Ni5x1Ec4Xb+JtNL3/9QovVP8N5j+/JrmwAcOvjSVhAyEDwgRcP/5FNbWxzctNpFVK
KIb414aWaCGUQCAStpWqFdpK317tD+RJ1z6g3cXQGmk97z4Ggd4n8DGKkAOAiU4jkzgiQWgCkBa7
BJSyvuej/OSUIEkZOBeSf6kbmfXfIBRDz0UNW4T1Cgd08rjx6nC3wIAfARFJQBXZPsC3vT7CwdSd
oaDaqk2cBkRj4wqbH6p3nz0Xzl4JIvJ7DQTdb2zJ1hD7mroMc3iy/gmuwBFjB8ul+qwE8KRfzGn9
HlckZJ2IVK9/1SzvVNzSIc0aZUKGGBKp2/dr7vOUrTDeeQOy512IXOK23opT+p696SNdzfl9iQNY
2cDXXXqyIzEfTjOYmuAmGsRtwRCH5vgB6G/wFkV3UX6DM018b4lLXFj6wtzUXDGutbgdY98oN5ty
uxmCcSSO3EF4uxYaHvWHipykd3la8D0VyQ8/gjKppdUQn/288EpIOLhy8dZPMaM9pZStlbJ+3TAM
OsDerDf41DXfwEI6V0aVRabJg3DufQW1XrnGgJ2oFmAOENlsf6oqE1bAENhA9aGlhkC5B4M+SsVA
h3ldIWT5fYaN2HetmcIWyrf8rvO29QuJvyzOWwMKrWN4qWl+hNIhTMRKyRJeKhe9Y/8l/v1r7G0a
+aXVMUoJRD/l+N/Kf0LtdZOmbO/8g4yLvVVBX05xUJeNMGhzg65cAw6gsde6JeBG85DDEkuuVY+a
Nub1h3gEt0/e1fE8+SbZBpri+KCN0I44SKmWm0I3wdN+xgck2UmM8ic5nP0Wttw2EowRPO2sFuvk
qFisSUoYV+xkRnqu6Hl4nIBC8BAe9IapmgPrUSxBWcbxobx48MGax4u0897+p1ik2oX8EsUex8il
4ZZs96DcYjAZVy+BiSL0+L0XynNHyFDw8zm8N3GFYDIed2jpiOebyGgb/ITFyX3m/HYyW6aayQ+p
6Igu4fx/Ynbquqg30fQeXw/rXPOPr+H9MMT89G4XC1e5+ANNVjBSrP+u7Oz3i5p0RpVdueI8pIrs
TPaGwce47NSgTPhYxEL5bs5Hzb0Z8Uh8tGd39TZnubaE+xxp7ibRCGjhsMMfDxWs6LiEPY1KRYAs
pIk/wORRoMaiLODpmuVXg9Dvg2pivS+m5eldMZbTCpLb+I9tSCgAiX0jkAqI7noWdUowJsJBw6+e
5M9qAWpw/yF38oKjnveR33EJJlhn56H0rhGB/9y6H+GkrpRgJhGnuAjpZYhbDjkf3ByS6C9ZxI2x
Q9bdlR7FPyfmVLNxTI6nNGtmicH4fQm2iIAl3e/ACheV7/S2AJ38guvDogKVr5RYf+joYAgHVPI/
xLpgT2xSB7VHSG1a0eZUiilr3aca64bvtyYQ4uwo35quqMT4nJiC9PM2pU6+0glHNHLAarnfBr3/
bijQkcG3jx+CEsm9I7B9LjR/JWEau5hPViPyDajrfhWn0JDriFfWRg2Na6GMzpCKY8NQ8fu6fWv3
xez5PwXvS0MpSj+c8mwIxcxJ8ANyJtMmsPH4H5R787zmnpD7ayB3viBGHa9a65yE2RJgmZZQjbti
ILaVSEy0W0v3SKcvyPwQnCP/zxS3qZVxEtgHSm1rVGVpgIhZ4GleYklYvH8RPTUak443oM7OQ9R8
Uf+Lb6P74/pBLleNUoIjW7BTJR8ag1Si+pmwCbpuuFvf7Cv00BWSyvPndMCifEd2sas+K59Xdt4w
vIK9TZU8v1b7S38GGK5MYzCuZE91pQ3VBR8c90mqALE7+O3/CMYxWZZkDMmp4ZjhaJsZbXdib5CU
50ZQzuoLIURXiQRLFPaBk7+t4/QQQezZgdFTL374N280XQwFNL1wjKQjXOuzQhIK7UQCCVsnBEht
j62BnRaxf+wm8s5v/E/TeTof4/YikFrFODG3oSYFWOjvjvFFgXQJSTyxKhsfgiQwIyHo8vroxEDz
nPPydNxD5TJIINXK5ZC9zjZf7z+BODhn4w+6xQSWot9c7FaE1tro3Y6pzNyqwcG7UByQdlqTb3Eq
JUQV/ahbMSRyr6oovU2KLkpe6ruQ6qAgC7CZPNRaBxZbLxRSSE+fDQuB13+eC7BPrUQZwUYSy9Rf
aRwC4ac46B+WoFsWCaZ1CMNisl1B9+TXe4O9lzOYQrdfzwHcAMFRv/rjPFGAkHjWs+G+X7lmFbD8
h/HkvjC1q+n3bNEzjfLmR/gxOR95FGEu8va4zavCMbwIjF12ZVJK5N2OckDu7BDRORHyx1Z28VqA
rcHyvnH16PyWUGynm0VtzyGMFagKHPO21vhqXx3lwdLjRtSBCjzwgz5IZTJ4GkVWnb3uaKRVq7dx
enJdFu95K1ZC7K89KmkPT2tebYVOtYrUUPNuAT/yye/UB8p9YRNKmZQ4ONRWsDP+ZEigJuqDCvg4
caofaP+XSUsCPlJKUKhn1uvnQ25nNib8H//918fzwr/0ZMsP2q4LzRoRd9HATZqECxjx3YWuADfg
6dh9hR2CwWRKfBh3FKQIrugfQmwd1klOgIlme64Yb2B+Ei7pnzceeYt8NVBqxtKo95zntsXuEUpN
P9SQCEkmsR8m1ElhtyVinMo6eig8bZzSbyUOZaTMzBWknLEzwzFDUh6lkv4DajdtDFee/Yctv28M
8GTWo8KULxGHhGV58tQgub4Yi5ltSU6v3j5VarX+sMNRFXBs1lMQ725qR6cZrNeDZpl2eKa4AfDw
iBkW6dukp1bKN8N4no6YeLpc8vgM/rA07GEDxQfFGQ9UcjcI5IDHE/pBJONJj+60L1lXJbR0RPLC
d6f4nUDsSzoUnGv/sMM8vQrR919Bzw8GEKKnOxtXjUp3Vvm2gcYFPizWqmWMHD1ElFx6PahLE3LT
4Mz0EZgKv2BtTMASrJPzrMZU84C/0OdFOpFE/e6eZniWFs68RIhn7En0Umg6CSENwFcDDFJMZhxW
Ll4U3a36b9knAJG3JqSUOWkikW3bi6+V8XRWRZ6i8E4ThZz16JDqutm4naeF7SHLPmORAMG8q+Xz
yO06tZkq64fTSiokEWO9xFU1+6gZSg4iVBJHrL0ILreUtom0N+8XK2v5b7M4XufUJvFIHq64DFBA
uV+a/iCx3WscySRVUFNyKsmihlixHSvj+iHXGpTSL41khpZ7dLXW4a5mFTtkTeZaut4TG0MN5LWm
+42/SXEOBhvDvY5DKZjhZGF6pbOKLOoBqMVnuEoTIInuunJWW0heiiSbrSw1I631R5IBrMvb41Cu
hU/lUgVMY8Urra7tgPVRCzTfopi3EcLflYdRU8PjqphKD+IVi8Uis94FaK6eEe9mbbmfDNOUGYbl
CrYACKhS2HuIjC6c/VwpIUvlVQh+voX3jqYe3EXloAN9IcQk8INnonPVLOlZqS5kS6Xz35Qs+HGh
LaGBo6VWcDbEIGop3goM3S7/lB/I4y/dIEdgRvNEPWnTfrDa4kaIrS53fHoveVMIa9iXpOfGA6Gl
m+sXqC6WAWzFu4Ixho3DiOjgCNMZy/HbSA2UqC9PVaMBpp/hkP7CLT5gVKhIzGIAA9sg9kE6z6ZZ
JWBCVWpiX9TpZgaosOpH5XqTvuhixKpoUOaucEJvdx/m7N321F6L6Jcon1JjNlyRhSZ26RHz7+q3
/W1JNYAU++UExoJfM1T934+gfVKx2a1z1Hx4f4hwlDAqOx8dv9ZnttFfX6WdGpeoiLxUU4eFjL1z
oFOw+/I4ikNePl8mt1pM46xcM5xDzqKOM+NmGJBqmbHerhRAK1DRTb8XNQzIbWQvOkAkvLZKjjwv
viulHU5FhWeuWUGRhVbcsdTMkOh93FFTcQyDc+ZxRMy/yGRw9GYulDoVdbpzzC5idW1Afm5TfTEC
r2m6ArcSYStPkNSzWvJhzMEVXXBbLnrY6mL46DfI8QHYYbPQ5wgAweAHDSktN45loFHkormElHBO
XkYl9sZX9FlYgdqIK0t2mC64WUs1sgbx5oVwx6wv1c9XZtaSHA7kcQR2h+Pc0XsRCoJm552d1zcO
t7FzYnMRSfPz+NLy9ridKUULD5eq7xA8j8fPXXl6ilAGZAA/v3B8oDRJBrB6shbkPro0MJFrS/2I
QfbxMN+G2T2o3cD3819GBr7SB+D1EG8XWRnOhjWXZ9GWJl/g7cAmiwoFqyxu5mDhgS+IAQlaawBU
Ky1R5gVlKicASH2AY+ElebvxmQYw5Kftset80+hDnxCrY6/3MDTLUrwGoUg0BjuVCu9hHF4dBnUk
s2UD1Z6iyoGEjvJqGQYipswCT3w1eQIGN0pU2cIFKNCztcU1+e0KjDGoRD/0wXytP/kHn+fGJPaP
KGCCD9NTze1hIMuivhIJwINAajv6/YS5DVdzN56HdeanLDkUzdDoXeXcaDJ/qp+5Cg2Hc+wYwA/3
Gusb2hTTdV7gS5H5b20HOZgPN/V0+CBylMVwF9nw9kq757ncFM4TVRW2yH0dX5hkwTRBCCQuTEo6
7nH4MqGDPIfhgpFivuFjUgtaOyT0FfvurkE2uKZgZQ0L3R/WXZNZIMfcrfaI2q+gsCHqKOkZrS6M
sRYDjRsRRbZ9hv0N3kSzuCjWD1AG8ttxcd5gCmzqqr4B/MTyiFgCaD1AmmP+8RjnTTFKmxcA78Ej
Tltm78w6ts9cOrgXBjEy+jZm4YCvsd1AT5h106djo1SvetqWgs8T1Hqpw2p7u2k9aCsr9jgKB7Lp
EK30oNeCk+IeVyWoWcRA3hLbN+OA0jss5fqCvgubhd30K7pNWydd1RXotGG6G7zjzMsJDIDC/lNO
1WqUsTCSS/vYLOEO3VzXGpuVealWLgtPs1YajkwzVtv5xg1ibcGCdSimtYtbaNjavH5mpOGz2tp1
eBT0G147TPZvnhslxyItadpUW3D58+BLjXo9jk5b8ktGZAt/4hdhYhrE3Tn9Q3X9JKMzPuCi0AKk
jwCEdDb7SWYNqqMvuH+H04N/uF4gSKUJ4z7Oozfe0xJDXvtfL3jIeZTUjLcXhUrn5xQDi2gqJp9Y
WmQw7iUQd3rQ4LlkR9/LfrIy2rWhnZq5mV9H6p4uBRid3AJ1UCyqbfAgmV2NxviNCPhlmy8o/HrJ
mi207yOVR3Y9BNyzkToc6N5Bg1zU/Se7CMpYXKVjl8V+2i2s6kdCBsaW9c7hxR+PIy+I58VKkpi1
2DEHKlBD9YvoJjavc3NxzpnRme/AHp/3sWM/5RGso9jfj843izvMvq2gZDzYugHPQfaaPB35L8mU
erGyBscZlneCAFMLjLnY3CfJXfEhMYwWQCmH/KuYE15lezVI8UbGNC2MCbVIrmaSuFq/VoFickUL
GiX2bBm8BTvGRJhvcw7wCL0SBNvqoL/y/udZBPIwIWP3f+CvvhoAfgLg7lNlHXjpijWGsvEYCpir
bheygkvDu/66kQeQX46+k3KwEUktE2RZiPah33dghGRXs/LwqaZP7mEocQ+MOEmwIdrXHs7byn8X
+WuOxfzGPCR2v0uZoyhJZWOmPPqhX5fbkSVWqvbqphgycyj+y+ImRnNLEb8RZ1auSwOMmADuQSDn
n2Ba7VNFK3pFKFQQKn/aIzvk06pkLRr2eEnXRztCs7mjX2HfyVmGEwOdZXhMkPuqC4AVD/rvZt+Y
Cw1Tdvf7Hq9nuoKVKu+BfQ8fUJrFCeqmFkfXjyl/ob4WpVrWCddeFje12BfSn0zzC6nwRp1Evveq
n2rkoQ8mUrIVY5H89NzuU1cFztd2mv7JwUrH07FdbSoG/T9KcN4MqzNltI/vS9j8BVKX97dhVWby
ZxI4CW0tSYPPQr5pRsJ/Xfc4anYnDOxZX4/OX6rG558McRLBfELtPM6EKaUr3OPALKdOCAWGx41D
t8ghB4ZX6li1SHzyRndj9b8t0OJUR6L8wo0gZyJPcjwSnrnBr0nU3EuJqJn2Jj71fN178/Z3MiDK
q82abvDnLAY9ePcGw1hg/PjK2doMg7lXhLg6UnAQrbZS5alLHbU8XjZ0MNESYeHQzZLaKWawlL7L
oI8u1zVYePPgdZzzk/D5DyUEL/+U5rkJIEEqQAkF7isF3ky80bh76/XRLBYlDTkcPWgfCHIcUxIm
loejthRBqw6+g1dGfihxrS+CRQroL6YsIGwg+SlebWNZ15lFRVRNwpranaZzDnQaXY8UpoOWFVU+
YAUdCdBShqw7XQ4Vy9aUag17QKFenahhD/sj+wPxzsgFakPAl8A7bdmGMPhKy0pHKs7QI+2OCFer
ZHD1qtAw9RAIbc010UNIYreXvrwP1gRDJ9KpgsdxxQkh7bU5sjFyXl56N0gXfJsDRHp9En+6l4RB
UueUjbekgG5Lag2m7Swf3Lnq1wLeOpETK43bXM6walFRd6wncLLzUPm4tQPillm9Y0UrPcaLsOm4
tZ2hm8VJmbwFE3JDdyR87R1xOu0zF5iING1SP/uobKRWkESoEhTzaf33Y4hkcJAyeXfRPCneWJJm
ApllZIqK2+rmXq7yBlPmFvNcRNtgr2kzDiXqTz/5shgf/yPlpux8Rdho+9An5DXbvMMbkX+K3lQH
XcwQeZLknYB3b02jmUkD0KMDn2hcAmJo2CTG33nW070aZtl3xXdGPq6LiYFl+0YvhEfWgk6JbBlA
fhd44hymAixE8Y7Ox/ysqfM9KKY3DNO9ma5Sk0RhY6t61r2NkbSJEwAYfmRmLLnKT+gLjiH0E9z8
aOwYUcWT0KTxht8XKFG6gBCpFhXVzL0YFuAdC677vJ+GMFSNrkOHphOek+8oT8wT5PR4USwqQYoi
gzFs5Z5Az3067Q/kIIuTG2GRaPetx8CKoJhAq5qaA5oCWEgV82Kje343xlomUjfHEGl9V64bGSOt
Q5HQkv2BSyFBNNWRY4h/uLQN0fYuAptiuDzwrS5bg+QyilAZmkpx8f5qdkUfEf//kMj4XFcGKl1E
j0sQDubvXG/g6FL96+CNtz85EfYYLj/Zbkvsxsq/jItTcXzekY3g0hjKhlSSqFoioBoivnSXTdt/
3ZCOOjGALH8ewepJXXdaDoMMiHHddhJeu2J9L1HxV3CcIiWC9eYNv+e+ejl2KSlzwqJX2AROnTDJ
XIsgJ348lN5L23eJqssR7Sql6ogCC3FPRgdJUeJH9h7M9BWW34S4oI8/3zITDen6zCS8Kk/XxF00
YW4lOTnYNyz5pGqIwQLlwZLRuFXLPZi2uPWI9n0ulQBq0gP5c2vGV4G8ucuPjKLryLBHNzyafVsu
loQKCHxqm6jZXXMxUAlrdtaFyzQ6h4TZrxSp/8E+EBPu3GEpH5TDAFFeYPe7BiuMYV31QO1A53CV
CPT+ICntR+O/Kp+69/vl9HL3QEV087qq8leIG7IimyBNroIXVZAEKJWzwjHpWz4GPLsfVmTcHwYK
94LymKLOm1p0znRw050prTuwohof309Tql1LrlTmFVjCC0Gzgu325tDAHWstPSbekUEftDOjWggG
y9dvktQo0cAxWBX8Lr741ppFiLhD221bjM+crr0vu4Wz6KaYS0guO4eErGaCFCCE0CUTKd3mSfju
yufGs8JBiuAzOQ2WBGhGJb9bHwzoohB7oi3jRhn4mOYps81n3oV2/id2yoZfv1l1no6/H2+Pyyva
9NbfjLzK/Eoo0xgVd9+Iu+hY11c9M9brpnwwIBBYm/OkoIVUK8DIRMPoDh04XaO4NFRdb9lviBZu
0Ygo9OIYpDkl+IFypA3J3n6rcAIk3NXAjj8zqxtLR+m4mMw16EExsTItCZEdpgR5p424Z/YaMpGp
0VfHqcS9N2palanWNzahgIe0UyCL3ymag3cA0HlLmTvwNMH6VNh5/dkbcrr/wP7t7JzzW04P0ESe
Jt9d0O52VNce49x7tqyAOIJyq7yJSJ3jZRUSfHAisBYqsIGI4CxjQtAgVpAN3olbidAUMp8/HU8l
yeBcihpwKL/VbXNXmfMZd2icGAiesxAev9C6KjbbfsIzD8xl4Ou/K9+TJnTaiRlXnQdoNrmg3d3o
JQR6kfo39wy8bLBwq90Ppmx89HmxakAEedraZx9EMiu7dTxmvStmf5Uptz9xxhLCSeV/obG9OQxS
S3nd7R3hTCgHD3Qsuw+E5n1quzYM5b/APGkCtlvV9Bb71uNP1wztni1LAGMf2tFC4VSh2ZEOWMMx
f6mk0JUb7IXzzhIRYxptwFP+iDkDCZlAkO6bNY5XGpbwicYdEdH+uiYkwv8j/CVtMlrc7i8LHXHP
PD5VcquXSScGobE3ZfCjF+Q2oIuLEiXnN5RWUrDdg/vkvBfeYJNC48Z5hFvKYx8ES2+NEWm0Qm4A
PWSog4WJAuLcUvujYORMRh66po0H3OkUsjFLXJIUSpiHBDL5JxIRlGPtVwaBxVLJnO/U6TMyspn+
rfkQIC4vfrWFuJiPT0i6rWIc8AFM8PI9rSAPrSHlSnRJheshx03GfoMGOUmOy1P7N/oDXr3Gsg1x
/lKOCtRdF4AaUC4MRAuKCkqkvmJs8tydc+N2o+cQvo0KyUJ2KFKA8AVjRyHZWrS/lWsNGwvPdwmU
ekTUcFmH0xySVk3lv8Qg7iESjs9bq55E0f3eP4j9jaDVpo2duYSsMGnsL0jf9AQ3EwiFBUS27LXw
IM01QEc3ojNZuy1KTffTUwt1O0UDLn/83fMpMbRFrSqAjQAFjcqAm2dewktbfMsBaTZRbqkhp3gj
Fq8yB1ZF5DDJ7ee770pPlDsZoWl5C+3WtDkMWKtWtNBZ4Gy9SSEJpSsGnyvPn+aXEi7NFgtVV4Xp
zSnnPJgEOMO+alxM07UIaFmTHb5+RikSRMwJKI6oHR8Ulz3gBoXkFEpqtQWw8xFt2lz8E3OyzVOp
cEvoRZ8AJcO/l29MFA+EVfQ9ZdZXeafLWNVc9DRngCr+3jOANdtWLk65Nirb/aG3Ge5FxlSmqCr4
u5Z8WicYM6pQF0UKhq0EY9+z/VbnXQB8m4UjKfCmC4Xkl5Ek10VXWy3Iko+qMF+oXbgD+BcqqXHn
RnnuAsWO2ci9BahB/DfqTZ4z+cW/cJogc3Hdzkiq5nVfLxKVwhTjnj0ZHEpU5jQf4n2CZXWOqxB7
xWIxn2RS9Lx25QgEDq4Ak5pcKuQcfrGumf5MO0vmHP0Z4yH7EUOJkebNqDDJsO5eZwegheirZmSM
+ngJCCNAc/6wSOqAKO6pRe3ZicAiW/I+j9VbSfDJqdnDPtunzstzlIRFceKGKPkGezdR94YDQ9xz
HrLO6pRhh2wGj4JreoGI8HJtZ0T8sUSLecWAsdPcl2LW1fj9rHlZZ5O+4acuna+fPyAMsaUlAgA7
HPrUO+ojttqC4egfmTzG2QGMXOx3xqfZC/BSKn95T4AwfcvHzXhob0dQLPdR7EbmxeHU/0AJFFl5
y2gt3+Ea7sSvWy89H20wJHCphSM/mIKoUZXY8wlUxrpfVeHULjxQ44pZB83DjpVFq7Jv6EoGQGXh
IEtsus0yPUf9OKdHvMorhyitSFHY2QUFEpeYHHudU5gqtAViImHT6+WDw5Sje4mYKylG9yGGm5V6
fX2VkuKzZi9Y42Nv+chRSurmD0PhXLAfysLwFNXXiX89/NvkB/W4JCk3QPIAdxU3a46p7srfdMqt
KpN8ltlFu34fAjSsSiWbgxt7qZbZECoVmQ+AlbyTYHrpfpzT1FNFVDF+aACfNcOqRyUnpLrrnZz1
CDql93OqUJsTxwDI/ih42uKO3aDMOQy7+N5SKi2TDfhNwgLtzAB6lXDupi3xlzdQVV7n58HfMgUy
FjcJB8QQ4NA9ka+wJuqYrH8QLIV9UiaURlGJuGRXKKR9JoqRaRzDOGmqZ666KXGUcX8lrPeSce8j
QsNtCpDWQzjJJA9pD65MDta2EOnXFyockmS4ByIr1Uc0+NUjY+ePhXNOmBBZQYv22o5CVwD0pUK3
J+CZka7WqexsczaSDm9jJb/tgy+PfVmDtRMYHktrQheufVXd8kVk1fmMgdpXS2B9b2d6bEZlDxYc
P2NvI5Y4tZvVxZiCc3u8CsPqfr3eJZzXtxzFmA5HoeDXpYy8v7Fxqc4kCNZJ8zyxrRxtbl3I/5Bm
5XlNxfmZNhZCihyr93hnb03k1pAF+SHP3YuR7gQ5hiOk48xwnit8uxzo5QxTuGKYUZzwtSS1qw8U
qYj7qB+u4pbxJk4uD9QywvWpgBIDMkOYgWJBiatKpobT262FMhTnL0wtQ97sixMVFwUf1h75vnT7
rT2nFjctELpf6pq9Us5dccdtue1omkBIoYsOHvv/9XQKvhLJOUyRXCdRR48giKxZQNuBejqhRiL2
BzTwczVVXfzBezVJbpFZmsyJlO7lPpoiq+mE+iVQtC6fkpKbcUZusHRRET56UJMr2UyfG8Ml1v4v
Hsu94p2lV55A4XF8mtVI7ei47pIPf3/RJIcu530PZld5dm1HhqjPn7Ifg/lXpqNKJ7ycQ65uwfWk
YTKDQWj6F6RbEZvNHY4AYs+8JBD0Da/naS/EysSVsCOzPukNVTJs8Xo+R2LYle++jvy4EQ1lYMJH
Xv+2FkchGryOT8jEVtx1MTpMJaHkXZugdgjH9EYEExos18Zb0E8CIsRRgx3h1FuRwZLGCUhidXrp
TN8tO/POEjc/jI0elkieHUeVDFiLD6cSwiuQLwZlmPcdNv5U2AzMm1NzJdHMK7TugbVzAIvl3o6d
wx/QDsJ/YayD4xf6yPzITm0eTgGKVUObnygbx8f7QCNT6ewtRihXODQ4cs7hnSt3Ow9lO4E2Y8F8
Ng6nL28NLrjAIW0LxUZemVnOuAIY1DU19SdbImVD8KW7II5TOk1ErtLSSxUqYOe6TSPwKJMFy8fd
djaWqU1rwDLnxx7qc/ougr9MswxpnpeFuMEwRHMGr3pXLb5zYNHgvOvgv1bOR3oiMxHsLzQv7JXa
wVT/6Ra9iP/vY2K8OwtMkfTx6tFcezVJWS6nbJjABMFGKjKypS1sksdBN5L2jM47G42AHD6y6R9c
6ePuJ20Dr2zsGDf22usgBr01Enq7Bt3uPFjENk0KIXCWOjXS9NuD3Dt/YULh2CikVvUaZTXBE76w
AgH7BoGwsxUHaa7j1FWtJxe5vExKv69ZbjnbMyYoXOpsvzk7ahHbinO3wTPz+HIq6iV99EW+Q48h
7NBoVLFfl7SXoFA3i8MAz3vi9Beir16fnqLD+hCUMb7FkuXFD7/AcJ4T9GD+l8I8Tt5kPYUkGMy4
qp72OEDayVoBdJ4uRjCmy67vXpxVLpNsJDES1IAS7nbvoM7vwGuiX9mdn/fjRzc4xxaCEaK32B+M
anWzNtcbTlrsSwDWTMYEb01AFafa7op/MhJfc98lwfZql75lJJbC/C/68wPeqgb3KNrypQ+wNBfp
FXofAEkMk3HStG/I/4OoXjviIH+q+RD/pq4Fxx62BaiikB8BTkEdAsxVtp9E7mdh4Idw/MvSkxEK
lmK2Dhdjtq1Cz4DHTR6VP3HwyjKBdVqNggBQ87sGDXmbvbwQcQeIQZvfu/2GYhxVjXvi28N6O+M3
WYsvS/fKu1BokoMIXvcMVXR3T98eBO1jdkCWXhyAVLyg0vV8kVh36xJAdk3UoMsuzQiidqkLQ5q1
ybAVDVVvn/vyxqEXdCDkRHyQJLcx1TjVA/DYR/M2iyKlQlvDi4Yjy/asuCAdcw2jzHIkT0LaqVEL
J5NL+RO6ZXws05okw1FZ4dpPKCIQDbAjzW6bgA87WUbGzju2U9Rz41qBc23dHlAMM+S1hqeoVCYd
u8Bl9iqkciWA5Rt5vH+4QhDkg+1eSTR70NlMhJX7S+0QhhGcVexU3IqU1cHWBDQoojbGkNVtbJLB
+i6losUKBhkhyxipAzGGY2SQdIthLlJ+hWmxx4yF/t1YtFlnkr+4SPSpv6+p+iatXts/0JLJ0Gyx
fygkE6eOcRj/SPg/CXhV8bUOVaJHN06bwgI4t+uCjKD8Nf5SHWo+dLVb8iVSGFjVGaPDZuJTSu1j
sqHZCkM9nOiutgGxHd/gxNPGYMgRamwHx6dGol3TYLdrDzo01SKMTB3X/baInQSeq15L++DBQUxk
/lXwYRZiBc57d6e1DYXfK2eFz1tDQlCWqV8zO4ErytvRCdempT9F5G6jctOTzDM2WEcfgLC0NTkd
mIUcHBC7Q7PChB8Um5PWxjgps3j6GASJapRWxeswRiZwK+cQOj/vAn2tDwlHal5cnvgbWRIcPbag
iiMX3Rb+2qZeWhJdlCaqdzXDOR1jLm1NCYLssoPv2DeZCljqftIUKSltPu2imsCy4WSGHFTae+H4
/NHOKkyH94zhmpyG55bbVyEHt+VvaGRIoJbg+4PUCS96I8yeQsj0yrwqyVj0ESi2qXsyNFMOpjm6
/XHfMe7ZMDcCMOOkS6YhXThDlRGlNmF/7ydmRhyTPNR9VMlzhh7HNsfnj2p93ggamJZk8of4ErPD
EiomPb7mkjedzeNZ274ls4kDm+EE7OLZB0fZ4VHEq86/NNs/JVIxdWL8/0cXPQBlDfmyOak+7CJp
22PViSp176YaiwK+8Vm16d5M+jHvu2BePUIhriqoq78O2ml4iJ2oF4BXff/qdI/gRozi+///8zRx
ich0JkZ89/4l0HvUmtXgraMY8yx+LDG5eCqFBqGhKjubAMBcbCeh/cpWnUxpe1gjdeN/YK+4QUlD
cwUktjTX9wbvomkDiEOXcIRcQvSeglDK5Hph576nzoRCAc6CAvO/wLCI2Q38JmWq4C8MrWX6RAMt
m8gcB6kbF8bP0hrst3zfUJeESLwQjFXq1yY2hZH286ngVxSADHb6Hq6dn22B4M9zSlRUaBSBVOFo
1+zTTJfEYTHaAzp4JCYDddKc4Ge7VmibHHzoBHgHNDYznIxIWsPVkrvkAneoQ+LTK/t4WeOaIv2Q
7YiU09mt/L4mowiRco226YNDT1EpHfjMwrDr7V1Q4q7ac9pbteUlXaOJUVj/YXcCjPAm6w0lOJvi
FvetQd8+WhC0S3g1CBasXHyYt5jjZNimt42mQG5LBpsC8jV5NcqHDQcjeXDJ3zzf/27b6xF6HCXv
OnNLmthKW8/lLRX9wKw9ISmm5B4kGqXnblWHi6IQ4T+hQsXH3kfJ3NCiOTJDMkzKBq+89THeduF2
q8UkB+zPmEx1gH8+RUAt4lg+zmnd+G0kOnNXGF6Tu9cc52MAAasUb1P8gyYSKF1NeQ/sYOD0LtAP
64Od55osNGizTTBDeXmpiQ93g1xbh6cBXaajkCdcnoj8QwO4pOZNCvtfYDOdAea5IBivKVUlPCCu
NVD5Tfudwpv5UFStn3RhSl3xhCjtm3w4BDqKoYlQNYkJji1oB9nCDU3KoKaSS263EJ9htV5jJty+
5iEcZL/fjf/SAkXSY0FBk+6AfioW34PooqjGVFdpZDgbUv3vg7j1773n+1MXuCfgEWgQpt//ev+R
fAvY8D0+Yu4iS0WKlzCDJbluBPN6u1QegJkSTX+ZWKuXVFgcr1So4FPmQ17JMIeEd35StRSYcAqA
+cl46sAXEajEa2vHx98re0IwetGwBm5Q0RdKzjhlSu7L6YrSQHDbfApyowO07IxHkA1bvgp/Rnc0
sXrIn9x4COmqmYeYkb+VaL8wi4BOt+smmprZ+wuzgbiWLxey5sCHnQYaj6W97q1U2cheBlRXKQ6v
GMldi2xK2myjgMFJEnH/9NkxQy+UP2fMc3RaE2V6lCfOskdFfCcNsO3kOBCMM2SrOYC8m8CATAcq
SFEDvsgtEBl4AEg82BeIg3oLz5xH+W9V939btD6u0ttCBWjysz969UJcidciEO7O2cIk6UT7LS61
epnWY0bCz6WOSaaD9MCG+78f/rfFVK1UhGvmMWDMZMTem5uGpNH9TUdLFCrGDARFhU5amSA6DfZI
5B9+Z+WYwnz3gNzyN3jSIMpemj+B7l3VwisCHius64TMZYFBdUQzIUgkp3z+nrOF8peIkEfjX2t+
02DZhsRz9eT3I531bUrQJIHOI39gE+xIs4nBJ2wSf1agQ4LxLyREg7l7v3DTZ8Od0T0+tWFkp3U+
g8/yg7LktTch3fwO+rRjRKahbuRpi62TdLqeGVieu1IxHWnwj+cefWb1yZAyU6rPBpPbQH3IY/A0
mtw0fNU1XdOhz6Bxyc1cyTSvaIjwWr6XqyTOkH7GwW2bQagujk9BpjdyEypzlLJj1cN2iHCHBmfO
lHD7Dl5cefOP1zGzb0lTX/z7ivTneQNy8I9x2hATyEdt6X6RSdDlLIBcgzyT7XyjdtulBB+QSOpj
F4WdMStCSByTi1Tr5YOKdTR90QWxZw88uHKSi3BtrK5mglbbRZ1GUpZcUDLJ5CRp+2DbMu6Pes73
I2f2vwAaKqva/SHsaaJsU9G9jl31FhHdJZbzJSmhCbPbOB8098Je2aGgT7XKzEMzwE93yTlzLXiC
3BJDZN8OSI/IyBnemuiABw2QKDa5GpnEv6/Tu68m08jRqaPwd/a8LuGv70vOo1SepNvul4PDj+qh
qikb0sDISZ+BxMWv02595r1pKw2v+ZXKKeJwJaUONq1xufifL06RPZnPSGwEBMjOQJXhPqheBcuN
2WOa8jHLdoRuMZknDIRxgfKAS1g+db4Yu0nwADOfXf0tdNwCM0XBUJd36uVhwIetKeBRQnFSX4P9
h+R3/iUWjfhCnssD/knY5kK6zLIUiVm9OFHbImpzhJiLbZX3XVxmVCpt1zh71/AjLx2I+3Nlubkk
MR53UL1dqdqf1xJ1zYfWSGVnF8pilw4ti76Jzkj5VMitRo4HseSLFsDWskxqm/uOUuBwMa4lggCt
WLPwtHOV+7y6Vwi5pwzetU3MqogxJVcEElJ1SXOcUcZ+wGJYblUKBsvFEkyjS2mVxA8d/F0GT1Lt
Xpi/XgO9odw/F30ZYjGEM9jbHWDSIEVco/P50pHWQXHzKpNjKPpPRaRgSHqnICX6FGp48aQult78
8sheDR2llIzV+sRzg7pNCdW3kpf6b1h1oKJuMS1J5VMJXt8+gM6CqRs/IH1vgvoSvXM56+WCJIa1
Lw1MQLxp7h0b8/lM6TaSzuXnf4bZVY60zkm2A/hN9sOa89PWsZc5bT4NJRJQoSw41PkloedG1ABF
eBn4FFKvQ82h7kXHb90C/8ala4ygwR2SWgvA6mfBkjGrAPVffDYnABdc53LpWvWAr+y5gWnBxeEN
qoaMR2BEIQqB8+oscOpDHGYTsPi2PyO5FZ5vIKzNwZFU30aiSvaVBJqkwYygk8Sann/ARAwegkoJ
iEP8Hp6pR0jINYkbNKzGD1RiTuXYHXrXSLHLVwgNk8q14foZoCCbv4GkjAxoWgLbwe2RmJXzkIW0
u71BQgamKOw8NIBK0GrgFadltaPz28dKtsuqlo7vNPx7yJkZeoInBYSYc2vGztt0YcPnT2MzX4qD
l1chYvKePDxotjhhOLQwjgJJPBfPdCxJmXYNknsW6mAhf+rrlU6XRXoDELMhZQZVvFfTLXKTtj18
aiCNBfafzLh7sz0WBddYGipZoxdVSbFXGVSFBDJQYx/kLHhRLxZ0CM6WnFiqgBDzLfaa6sSbGKZ4
2qmVivL6WkNTjNXuvGcFRC8qJBfrkj7TQ/5QW5Gue/1ySfD1oB+dbjJD+9GjrCWqWRp91cSTPFXf
g9lLVQ5dqqonqGW+DaHxkaEXFoAzlgD4ca+oh+YYgBmcyvgYfg1jML6XRbeWBRUbQBwXqKUgT4Xy
KJJbKa1SCLPAo9YAkooq/PeqYhpPwDrXB4SE0JH9QSEkyYtOb+JKPt+GbOfedXaiSWsP6hAXoxEZ
dPTC0hLNz2CDkSdf+SqWVGt5n7wKou+o0/rfYbttV/okzPlaSYSim240kCB8Q9dPiS3dVjpNg+OW
UDNvRcr4Pkt6Vj6uBwYWrK9I4hu2y9wjaD0lzDJQ/pE08aMxgaSTTHs80miLa1Mvl0eq/I0gWUlP
htKhhmR3mjuzIdliQofDIdQpYLGhc0Msjk/Hw3oX6MYYZQL4ZoWJ1W0ZCodITbwmJN2ZAX6SyvQF
kHn/ZmQH9S8flOKIjwISzPFh/QIKbgzMk5VbQ5iFedyqTmqtfz6SQveBeXWxYrZIUURodg5z8AiY
/kppjqeKo1uhWgP5I1Mt1qIKfxF/9+cf1oBAGPdJBB0ofDRhvSxVrCoOamjBHR1xPBzkz2G+H/tQ
SFXSTr+pw7je7DLiNKq2Udmh4jlW+E99WbwsU3Dbs+AUHEfocXgqoEzbJbAGuulPE9X2z0q9oOsw
8C8tQHdDRx6hWYrBT68F31CfE8OYsuIl9PjN/5gZMGN7C4cNvb5NwfyYHlJJA89j+WwlpqZtq+nh
l261qXevXEiHRxrrJUIhcWB+glTxAPxGpnNxpGGzxzi5MSRxdgkPNy7V4GHFhatQt3kGkKfMcfdS
AsRjZnVIY1vs0fqWdOjObJvJb+MrVZgfl53dYHWfqBQeAWulBN5JcZ6gKCVkV12qdUkRVJ5Z7Zvg
afHNg35FrNJ0Ecs/+E4VbZBJqKkMeO7oiG12w8rd250ah5WqotJw/edZudwZ1By3mvL5lLjChWDK
gj/5xzd0jBPAr6f/kOERnm9mq1kn5GsHxu6v2rhr36U0/wZ5yJnc7DTtjGP66NjtVPmirCiLJJFm
ASFMNIB2/Mm+InmRe0It76dFq6xphMyaDOUKURvUrpTgL9/O10T+Y41LZ5M9pUBWcID5GiI0riH3
sKgIpkOXknRcWDhdA89/LWtEybnzzyXF85gm8dShvh2b4vZ+YIfSr+TFCYURykm2TTYkdbOfO5BD
KEiyFO6V8UUs/XGZgij+akwahrthOzGhg8XLP7N4DSMhJwKgH48C+HRT9A3V0Kthkk8FLrS+t18z
TL3AQZo9gPkeWSdaoYeygjXK41FXvT90la5pddyYXUy5k+3KdKvfEEoBavWA4A2pvRWWcU11mKdi
5Vj/YJTJv6TxiwGxv9UhT2A99p7nZYsrNilRIJDbXS/LXcqGeyjUCkyW3qaM1ewxr/oSIkYCHnf8
f40PsbxO3mm4zJcIn7oX9oDWb3lzGpRfpyMXBL6ideJqa5wunkEHKrUXk2S2kYIphPYTvGjMY56i
sr+r2XeGcRgK/SecY3BxQKiJxCrzeqPda+d/5T7jYMu1S6pTglmKazdNvMb8qW5mMXLwKkyGtym2
JS/4qwzsBuQehcOBjlwFt4hp9M7SfrfoyxBmpe+wlmQJeHio/tiXnWIDcUMZUhEOq60wv9/sxVQm
SakzxHP3ubriMqejPvRtW/tDwkzYmPJQJUjsHIuST4iIEAKx6Y4TiM/zaHFYO5tQ4HJBinivk1ad
4X2RBQ2vr6carCg1uezOkmWyDE1k8NdI7MoVrDwwgr+r9wPzoqQBg5DrlTG8U0uvlDd00S3qEHYX
pPxoDVFb2QXNCiEaLPP5qux6BmHrMnMcjyziOL8/TB1qGcm4TIuau3ARSayxJH555QiwrrUN5KPd
RIE6dNyKLiD5z1mtA1aK1Nm1SXGh0MsGU8QwSZuLzxM+AUnzQ7Rf8NJgwZyP8TkdDhGnQ7SPCnmk
TeISr1sVlSPpA80JTGzr15171IZvSA796RXv2IdgVSJ2OdjzZtVYZtXh2WrUziaeGN8dvauH0r7Q
c9gWodgB7HTfGlbtRxSMaPsmZ8bY0qtWP9esc9iqvOF62bMyUUafydnkr4peurh/dPMHxUqd3Tk0
msv8xEa7gnmeSOMmEBIoyxPMg6OqH8atgNPznMV2VSJoR4fcaSqWvMuY5sF5vpO7gXRW3l/MHfxm
I8768gdaiiph9+2MyEE4Wrw4k8zsq6fhn8C0MvDK9uDjxmcQjIpSfnpXXkrP4HBzEeeI1QxMECOj
8OCS/7jmOIDbiCPnZtWowMva39ST/GVR7m333FPqCYS/rkUJM0rxSPJZJK7PmI8rH2+WVLNPfdV/
BUoqiHMbWbL2lUFDvvNK+2pTsjsWnnecCoo7MUyAtJtWYEWz/wIXrj1XhUzjBdhqdsX+BP7JPqew
GljoG6wC4t4ITZmeAxsCDLBr5NIlhannbm/7QZgVTCvzfCnqciUmfaC7+RynITHtpAe6jrxgXdYP
pEzke89Y28jJMRzZ1TKSAhOxKxTxJaga6gy6p4wNRYOLJr2ZIjYL2AyM5b6nlxRWUBSYwfLKaU0q
PsaZxAaSA0EgGnKUB2akkcdrNod/qMN5SBoUkA/HtXOOqk+hCZrnxOysUfTS7Xp64f32dP97qaG6
/rhzOjn6qgGs6diluH9+Ef/MLixK+cTC4iKSoIDR5kh7MEeUtB63LvP9M8oP9izRYywpMIzpzZt2
tbi4WLGBLnsdqnABAuHgCy0EqvTZ8DpHuo6xDTV5rDiSxrWi4axGNcCzXaK3cKeAyVXzHrxXxG9w
ICZzaEUxXc7qAm1b1Ocjp+BKCu3K63oEBppm7lkd2kX8IqCbv0ZwckQDrEfeI06Q0tLKRcs+bLNV
FFcN92En9iiXecsD1dO6AkMmaOQEpXizPZ3SJZXoOjRP1E2eOisdngkVooh97cK0zNITn8cN+pFE
TXy07ot1FPZcN76HSOMnCSxl39b5W3MF32c/PabxQTX7f+cWhy6S+6Nk6iaZewth5rTshFcmKeO0
mjZ251Fhu8i8DCzvIcfQq0lPZURGCWOUqnUnxFmjAfpRzmSZ17RBp2syIdCfuK6LFzWm8xNqxwGo
Vq9JJRVoNVUhuSrBH4DkytRAjfvCPu975q/4jz0wD3hfP3g3G2mZtw46LZtUpdQq4pvDNI7bK5KP
oOebCs50PG2oZ//uZuYjNZqK0Eyjo5k+Vv6Hpbieot+0RRnCVLH8rKbPy8VoZcEJihgu2tyZZem0
fUqSrOmk1g18dj9O8c6NqfHb5KpLmT/Lji1xMYs+TFe6lrBEBnyk0Zg4iFb1QZuNB+z7npIr2e71
QGrNJFMVhHbpeB/2Y/BIqJpr7P/7HRPsUIeSIxFLh7m5n/QWWAthsrRx1v73EeS2bs65QZeVRsRt
JVPmZ6gW3rheOp625mMRrimltuDOiOcKAhtOaqCKKhx62ajJ6e77t0RerV3oaqMixgPa/G7UtQbd
G/jiTPCI9M3CVk8M2rNqfw2cYWhvlISE0khR2zegHvmKBoR/Y2eEhtqwxnnjtg90wIJPjqk0MuJa
b42pgm8LRvM7IapV8eV3xb/arMCBf6OpNM225dWAnId/VXeP0jNMkbAJNWe4ubGOQv82hDJpIUbZ
KPlsQrZC2XLSAjxg0Q1FaSw5LIWWpxab3NqoOlujjPqC42+aoEozQ47/BGKaULyZzVr+JMpIoxY8
IsonKH7+JYW4BF2Eot1adlGkqHeV2o1QWbf9R3TaBD4DdDS9jD5wOVwCub3t3qooiLiPJlXHXxlh
Cdxi+aVQnv7mXwYDmu7Mv0zemo3Ntrp7tUwkD1BjhNYVT1HskNJFr7HAbWoiKY5n4kOJuBIZ1WZo
2XKwxofH6IhHg26VvKmbZcetf9tBjwp60oJD1Fcj0ZUMjOlax9/308+9lEMLfjRXPCbwnresfoq/
WFS0VIBIBlS3mAoPEsZxuhm++YihF5NLDzxxTsGePmQ/is1Lc7pRTkM8IeN5E3Nt3riiFz8pXLpA
2YK57gI70vvuKzlO8ZjQ2YMxB1RicWbx78HdTLqEIYX8XVFK05qDmKFqA7Y+Plv6MYKzUiLEH7fA
CaxcNjZ7odJ0+6dykNCmJ5aFm7zyg1PIzGyPprNbIEuFjr+3zSESIizJDXvnEdT/ggVFH8IL1z1W
DrIG8mCZ2fuyPRH7RylILmF06QuMgUxujDIy2jLU1H7o8l8LLh/imbU3jQxFHBLXXcJjduVmGiSs
UbMaQY9zCgWE8l/KlwlCzMIGh4gFjlC3vbp5oudsCCX5xAZPQNaxcp8QS0W/GLVFKSRLgN43Wtne
5aUEhlfO09kCh0MkmjqIVnd7PoIiSVh6ePsv36LYmRnsQKo0AIwDv+WYXBs/MctWfaG46iYWcFUN
Rfgnabs9uSwPEnP0TrTAj0RhgJ2aamCNuIZ7wD8Dqnv/gUiB/HLgHaBogO9p22LUwHvee91tDrxY
JF5SMmFQ7DX6WUv6juWv2WX6R8RBw3pX5L967CDqaYkVagMQpOaeU2n4Cb5O0OYj5F7NEWvgqj33
H7z6HVUQ6WNck0qWDStTzrCwqk2wkU4Pwtd1sszuj3EUOm0Uc9WWsMiMJ7aV/Af1QxdsSfxA42fT
0NihPd3bg1tNnnDE/Gbg4OtOkvbt55q3zu2FUtYawNBZcZplZPH9dHPJhuJYaTSPnJSQcRA2FSrn
KzEHas9gTY1is1Ag9cp4JJyDVJ396TrzrXwqe2NX6xOdF/qF7fQArt28tjKARR+Z5arf/KaHdkis
o7NlkjJitazDeXNwsfpUFqOCiY9PpwhDsvKI1kUtr3ADec0nki68LWdqHeFK6ZPrdM2XxC0wij8g
SivKttU1iP/vlqj5sfGLizOnPE+g1nOiJgFyrXdA3t6wCRq8KmgBLCIfy5G75NwfjlPz7kcRDfTH
ubstlv+MhItU1mQS8eeVXl3EdUAKdifselM4aocdLxjSr6qNdyBFEJO3lSp+nlqajDn76n8UJfMe
B+976O2rG1HXE+8OyIycFYusHgEvzVJ+nDjOAJhlsSlV3pRV8sN1SAH7O1yN10sp9b9X6OJOieIB
WCSmecsha7M7rrUwSkv8CX1iDfBoJ4ZNbU17nITeZdx7eIPtKo3lg+rC6XBjKvEN1+bKAq3WPN4p
deQgvnHHvQoQcYRLYLHnlY0VKnoVYpALZfHDF9vj3D0tqEBHvJkJBQQ5lGXtX5lGF9y4cUlyx6M8
om6qP5WSA5QfeGPKtPwuQj3jOOsWzqHCoI3LbZvCFouRgfUQeJTPqIgYgIr1YWvXw5K2KW0rggxp
6DE/39FrIwiUjam7PHghxa86AHkhMyEz4Uui/s7pCyPBKfgiM1lidlALhI+JPn/l7BTZpEvzLd+F
NPZYvzpSyeQK1n31Y0JSquSGFD/xZ8qVQAopJDY2rXFAf8VFNzv+IJVaVgqJZ9eQ2Wkq7YH5+oD9
MFz+QWgFq6GWxR/O6x1u3zLs5oK30rIC3AW2g5eA/y2y5Jr5sSshIBxcJbwO0nNv6nvoazFfcqtK
x7FtOQI/TTWfcxRSyrT1xpnUHe5nBz0+ENKuUvuOdZIuQ77g7ZqAOHxPEAaN50039CbE8VksvQBx
0f2NYop7/4gsiA3ppe4Rq+R6BOS0XxBp/SPh3/ar/M6U7UqIyJCUuHvXiEedDlchEezvAnMNRhN7
xUzCnxgzpgkIhhFUvQhVb9z021jOaoEm3pUayBSBLHtgxDyfnmzQtUZLgmwRX5TwvU2MkqzcxfdX
jopkylccLgrGVQHPTxn91KSb6wJ2/UNJR4Fp1DI++VMofFI72qUveY6DYQdTeadRWvmtUGsGryhp
tZdsREDHH7wHsq1w6LLf+TZOurHrsvbf5Lds2FbX5Ulb5KkuBsaU4A5ex4BJKau78jX90IQb+Teb
1PXztw/jEA6yvq9OS7cqBffM3LyeuE3RkR0qDiyDNoWQFcYohmUSpn+Vshkezw9EeQyfNV2YoqVc
1RpIiRgJ7oOjJcBr94p8cDwJJYLKPPaEZJNytcvd03XyIwi/23a8HIyf5TEzqGo430tdg/tH5s7w
nj3o5SYVIKW5U6H7/ETK5drqPA9TELFysoa9s3OQbA7qnAXaUHHHb1Vcf81keXWMOWxMAxBUR60g
diFbgFLMv0aetK1Un1swTssQYkFWd6ToM5PRKM41XQjKA493260ejcEcNgGAqs4E6vcQWRYlqLdu
bJiKNVqD/M5vDgVHimQLKQy+foUsCWs9CMrDWwNYZDzKsFUWUFlF2SdqOAI6NlWbtrxPFJQpwbTm
3KW+kSZtsvPMhHJvUSqKz6Il2E37tEGrZ+yf+0o83lb990kLfZ4B38m77UJyF0Qtcz6P1a9HKY10
nrokF5Zbkj1MIHVWreZ+7EzYXqnDAGytURRQIyLLFWvi4BOEyQO+cGH+1p2N0HC5nFoad76lmjxy
Q3tdhpEZGgcrG1sp5uIhGjplM3wXn/PDf2TwgX6OgnxG86RL4TYW+Mf5Ju26NaC7NPc8kJPJvC7P
Dlv0ZBh2/4pCmOIe64o63UboHv6f1EP+YntQEqAhEdxgN6AFU30YsCDCIC63fLb91MVCJqMztFO2
75LVxt72dzGDxTUAC0V0RHCTD+citaYbN9N8PCtFAcNwx760Cp9l+NePlmqtNEb2BXOvXGpWdi+U
mByLi3mEvE/XK6CiU1IOWEzgUR56LIyi9thbAVbnujrFfg1LpkPF+yfjlUJYjl+aeVmqTYeqHlal
ToC7BGcQ5tcdl1x3rALIMaJur0swLWcw35jKf/uYIHdsHLe67ZI55y1p3xQP/1QU6kI0C7naH4jU
pRFyRlHlsl6FoMNWc02XBsly7Xy0WtyBrjE2Y5j/r6EAQvwIoteUkCmvTjOssUqD2VJ15gD9IQvO
Gmlhnr0/TyTVGx4zklQ1iseLNopTcn73LvDIz5flGGJxyjsDWjy0D2byhzKoAHbGk/+/SxzWzQMN
u1T508L6CfQi9bYuLouLCaKE/khh5EgKjEHcQSAbDArOn9iuMlnjIhkzbfDZssTpEnPUOlBFPNmd
fo3y2SuOIhEqjkEpkPn5mDfV+OLekk9Jkg8Ho6T5+ZSJ/9XchbMK6qi6VJG8pD0ytC4Ya2krkECJ
xQealHdXwvCGBE7GI1p9onKfG4SJmtdWQZYMdo9sEjs6jWy9cLgO5vKWuiIx4mXjV8mz/vaBtyql
Sl6cJkmlVcIpwq1NjKHSMFwVcO3mkDwAK5Ji+jPhTpnUC8Bz1YdEs8/LYohD6OQ8GJYVDhgtEIAn
7ODcdOvC5bsDjdyOz7Lt+gbdlVZkojVpAyU/oUiuID4y6iytadfBazpjWd1X/GbgEaZmhZDxQlxH
IDdvdwihU0KO3HVgmmYhTtXhhvNc5ooa+HqdgXYRUu+PiYf/WPg66KYgDIkXknOVK7P+ce1oNPse
Qrils8HyD2eU+OfS2OatChxnH8xNWF+39cHmravBULs9SK4Uxzhauj+BscwkfnVPd5R9/LbseADu
cN8puSiYDRsh7jfLAvGr390Rjj4/8FSpJzcR19yhu1hs1nzErGd0v/4RN93n+ILVVXvauqlFtkEY
znAeEIAZKlOspP9JcEZDtjySK43BsxAhDKzdVJketFUdm/2n7xNbnbj76mkpBbTzmgY4illulPAE
k/QH+C71+GVfvXpz1Q5y9Bx92CS/Y8UYXG6yY1YOMXQRoCT/GLYicBXkbxwW6PLQvv890128u8vz
WtI9e4LzU9SIOPyQA8iH1g0qsKAS73T6P4hj+06J6KJfFZfE9CKGwpoQuqLYzbOyOyixw/3SJSV9
IhFFpkG/UvBAUHv/RLAcjLv283FwtnJ/bkJfdQyrhwaQC32nVf51SIsOsFCVPwgsO2NLH8IXfump
cN8YOpIIFjLl0m5bzR1t0sWljjjD1FTUNrrS/bIM8F8+ee3ZZOXa/2TgMpl1V+6keK5jG3oSeNGW
E7vX38RtUT3Zj0WO/gHYX3da3zRkpfeu/+pcD8rB7OB6o2v+p98459NCVJEOHYod/3Fsftc62gcM
zfhOtOa8O3XDt0sPEJA1Pd+e1k833jAs01cYaWgpCFJQwAOkw6w5Pz5o4E2E5k2qq4r4IKW/Pldh
zu8Bzv6gl0l6TgX/FoJfPPCbxpsn7vJfNwbWZ2mfE+6klEUdXmWV8RtLmtoX1dFeVj9dHdooIlsS
sQ4gIJ68URCUiPhRY8HLEGwZ8oAMxHApDCaAA6L9GfhL+3Ut29DkrR2w1UWe8x9wZS6aQA3tUthI
1U8qKEKsxs11U3ytcV6neHPF+h/dNoOp/ryhCbNvN0kbepoCI+4NJOJtQ3W4jZeiRYF2ersQgnLk
qB2L0u0t7I47Al07yV4JjoL1cOr7LLQvFexc71jzLbIS7hvrHLv2wsPPwig3+yICGaQqj1AOybd6
7nHFH/YbGP9wugjjjLYAdAJ8fk1WB3aAjrxwjKhhvK71EIBOiakrg84lySoLnbYTNJ4w6Fv9wQlY
+HjuukOl91c1ptScjqqZkPUVZ94IXCZIkN5DvhRT3Lw9hTxQAZCmLQZjuhvFtLKjPxlQv/LuNEb4
0/JgidbFbRVIeC1Hzn6s+81rgO1zi/uH6LG9I4ndrdA3La+kAc2VMbWzOZPx3I3ntdLBsN9xWpqJ
63TlKPdd3aD64Jh005E06yRJuVZxF/I1h+hPEjZvoMEmoK/rZbMEaDZtu5EM/aeSu+dE7xpT8YbO
ipuxRyXojDdoOmXNCB51KiT3RUxFMTIp214IWhm6qsZRWFfFmZbiRDCkrmdrbJLGysrBNe7F90gL
HnX9BYz0u6cQqIPSWpvPUtZT7hMVvOfzcoAR73tUYs95KW6Y9L1guy1W7Aj4aIf4vHOse/Pda2yb
6qif3qqOWTCC2dBUSNrOGPgaAUWc1NYRfEu6sRn4adWNZ5ZK6kmuj68SU9WNXSoql+z0Wo0Aqcpq
Id/3L4VxCNTAVH1dDBKlscWsxCO8hfsrsB2qLm+u5XBS7rYdwX46apld4twJBP5rKhGuHPl7rC89
rL5eopVNnDDXVS3YmLp5ZW3d+OssYF1qlxbnCvH6zwZ3YUNtodl1PyaKhkHzbWWKqYf+JJbB4q0R
+943nTrTtbOPaPTGgKkuy7am0z0HpaubLdo4vWBKPSaHnYqemPetToljZaR0CSyyb035B9l8dZ4r
lkChk6FLOYCD/gkovohGZJIwssevylcMqQs5D9tAvmCRDByFsQKbIP4lNIuydCrduXzZKdhIAg15
zhYOQ78CcKnpWARikDmbWAZnXpDOs1BoMY1VCxwjJ+axvNx8LPwbsr/d2uydDQGDnF4yIPlowFyR
8IcgTSnhKf7/3OzcgQZ00Ob9jlre/228UoWY7AKvltP+OTplk7nZC8bfzH//vUbGC9djyOWT0dpp
o9NzJL1XG1VsG69nL8uiW6I/XajpHeKXdQE7TA+Fd55pfOodeQk+Iwddzu3y1K6o25r3AeFe/kGQ
FBcPeodXBuBM6H+HmGzOePY7yZsR3Hnjl1MDlMJm1+U6SVZTbs+eSq7PIseSUsNgZGIGV8a3KK2e
EoZwTYSmHIW+7TUhhtJKiIfhbedfr3Iji2mbcsCHhbs9EHbuKax9gB0Ws5p2iR5vT+nuWAbiFqIA
OtbeZN0i6sgOS7Ns8TUhvDhzNLz7JvPNzL542WZRwzyc2ThEIuMFz1n5X8FzwK+WzaFxNyqWyEtp
q/BLIuVtdbfEnffUvOBUO6Ef1iSLmRXMOfNY20gww0ppYLqT79Oond4ZC+Uxv7PfEmKdcK3NwZUm
7sKQ/clU0DFLvDfFGF4nR1UHADZG94JP+ovaPfmRbgN28PvQZdD/n4raKO+kKJ4PM8DmwOd2aBL2
3myAKjkb0dT04JzfUuCcb3FDyM39+RsyLUIKEZPjrYk76EIdXC15N5sVFXoyt1kZDCJucmuzPY+E
iTf4fqj6KMzJNgTbyZ0n/2QwEC+BCH5MxrJOsdrMar3ObKY6amvKJbfFRvppTDO2NmUa+ElFkHOc
jnfKAXShZuewrmuyadOiBCmBB/966Wi1WQD40ADXRMx7Cdp4xOdTyKFp2sGvT4C5CV/ixC8jsNdz
KjFUnbjjU4xiRCCJBFtNcRdnnpS6l3V8X4er+Ti7u2pgGXOjK9LiTpYspmGwvCDJBSfA16SPC7M0
pFBoPCoN/+Gh936dzgBLInTcFUDpEucVq04klTw/4f7lxpfulUvr756nC7w8fxIXI4n5n+UJQFLL
dUp3yncyfJmIYDw47DYXEQM0wY6cMBxB1DI01xSn34QAcpzTceTeR6JKIkIO9BuBWRb7aqPPlvic
6TqziUPipd4FeZx6SiePLxrlZcRNxuY0iqYzF6+ftqjNbsAXTKIS+GrpmdQosJgk5SlOKEqP7Qko
K7ANrLBZETj9jSb7qlaelBW1pGg9u/NHqfLCDuhG3OfB+xGHis0D9uYFg90mGvfF2APR1xyveKB/
+bTrqPE89+7yGm2t1UezF26j5IYQOYXgwTkXjjwWdjZSq/rFLUVJoeqmyYpCu4Zfv5SU6RBSSyOq
JdR5eAbFXLL/lgC2RaPUdvTZ2o7U0kz2hfa61JaMYDQgtIqce28Rwribf9QRcocRRvnLucSnHb31
Usox0ifCp0CWS7NT0AEp6aZCMeA5UD5p0LJbUICBd6ErqV2oMjHp+f8aovOSd+33R3WDNNVo9lyI
sYPeWZAIrwE6xVZa+PGq0WSCJ3N6Zc+vgEEn3KNo+tftrJ1ppqIq+ye2z4VUX6WRhFHIyDelr+j1
TuaR636PpCQ0/MxUdWUGzixgNwypN6MwVVQJxUNzpN5BRGM0y1gZYzrMZOYEa1abpl30KVXmz/TP
2+kboSuUFO2Z61+BBEje1hY0HXeXJ4BMvIOaqZ26oM8SRiTYfW4cTDXrjmqbCEWtLwGhY112Sdaw
pakYU4QvGbOTY4yZXvlC+5JNJ/03pk3aihzBoVxcmFU0rv85uqW/2x0rOIj9Dx58E9G7+6y6w9U4
XJyBy1V7fRWElu5lcRYo/KVeWwi0mMBBd5GdumOaX35J0hMPP3VoinIrq0f95JPjYakwoN4K7FvC
KNI3h7iTB4FPnDo+8YpWcdcmH8KhSzKD8R7X957nV1mHpp4nhHK3Vf+akJJikVx5iCCRJ4sj0tSh
loOJLH6KnPwbUANmaWz6ZHFoXERQjxSLiUyjQF4to/VeArDBceSFLu/le6owIeLaZ5ZR7na+s1lc
Hnv4qMVP7T56b+748X5Su1AFevltXBbyqwXXILjqGOC1Geh7zAL3ZO0NuSzpccLl5FW+fJcYC3jq
PfsorClZV3v/mioP7PW7HdgzYQjrTwlph+lpHyWhvBvruw54V+u7KwF6mU9s62hI5Ps1KLEEMqcJ
2gITqoqgaX6/VknoOmebxUwUPf06mF1QRThoWh6ZkxNeHxp+zQjvCnxsh0SZCLaaj2XEstzN9FUD
Jjt+cMAv6TeqOT9A8gqxDJJBRoYoiFLINTnQuqAfIMhSVMEdf/E8jnG7Pua/pJTj6w2bP2wM0VM1
e5vLotdz+DuGnSXiyPEB7grvp4VS9W3OZExVWd7ocrKX7VT0FVfY7rBUkclpvSb2vsZ4mglEvKIF
70McqjtrYjUYekFlMXbeBeuWEhjZq9zDB6J5ErL0IxvOT4cLjth4Aqb8Eueuy1GWzYrP2wFVu5Dn
KQgupRIQRBgPU1aIquRLWFKBfBEOCwZLiFDFALpU+oWp2Ge39QiUPLQ4r/JLOEEIbkBD75livuwI
aOndL0L58f9GqzgxePxhGmb47P8GFWlnjiWQ/cHI1ELCVyv+YJKDsfjIfggyVREVndRwMZEdPAYn
8izKBJuzp5sGtBfmIZPgt9Qc6CtM45uxsQsjHhyH2WaEktGdozOH7ilzte+F0WWkJGjwuwoN1vrN
9YVFrnFf1q+kiLUt83ERGOt9NxMIHnGFpUYmU+0JrAkv/uKmrQqQ0iTNKvUYjH6LYuzlE6OeLxfM
dMdLJHdJjg7oz9Dx/GW2jIDDi3GEfLu0j6VkHfSzsngJ21WTA4xP2pOK8V5bF56gp1cp/5+QXUb6
qIbj2XJ6pdZU41wBfGxQLGeBUnfWH5NexKSeerNd4CfV8bcONZOgntqABPl7bdEW448pigvPfOzt
bqrp+/M3C3qlJ8Qq2i6cnzrjfS/CV85iXuL26d8j3XzoWII4ul4fczZsCefN4oLAIhvXARm14slM
PIRmqOJOzLac+YBuA/NWZDasunTQlCUQQcax6HK5ZstRBYYoNOPz8L0IfNtBp7AcsXwjRN6ADJA+
ayBk1S6+aud8v1uKfaLswlVsFPXZ1jRq94duMYddiG+AtVR/YtRiPcRIB25cvPsNcfjvWZSA8LW+
+hNGsY264m5X3qxdU0gL+w0GLBjKRdifjjWQNxZg5OPszhQ7BYsvSI1zOI3ItOGJG21qb4RD3OEC
KDyYgrZi21qkrHaFvqL/xfVulr0zSgYALFavdXZdw8JZHroszl9P5QI33Ax+2tpfRLvYHIf3JIUW
U6l141AQn/oGTYrDW8ZKonwpF2NGHr0qFAM6iZMw0w6tmg8jdkXJbjk4DP2LNeCkW2chxzipBixI
JKLnLAkZAKWPb7eHSCt07iRkdApnNBNnycjAnVJoDjEDO7a72gQUbL/+uS8e38P+H+Rrc+OTMEIz
VtedAcQkpg5RJATs83vG8cvhyRYeLVUWUWIoGWPz6Hrv/X4TPBG2QPzw6jU/zIo5lhugXwqJhMUT
rt8IlHNfKCsoylNr4sn6zvyxiFIrFysD9OwX8ib5zrEFYnTvT7JVVV2bXIFjiWvOcnmWjY7uPQ7j
V+Mf8A9ypTKkXlABgc793IvLaTNDcaoiAqDakwEkk3oV8b1H/dwl/WIsIpc0fwzWJ+Otro5gYTTo
aToH7nX9dCeyLcYEnOAXHVX9RH1csbb4qs/vH38+STTfPYbjEGeLwXOKRUy0Aif8KRIYXRwow3fB
0ZWbTGekzYPPy6qVazLi2rOmw9LPyw9hat8mdPcTMTEEj1i2x1lqxLcP5NdpppTVkVobIKFn4tHx
XNIalaNzXtpHgWRHUlx/ZAHqZd4QnAuoU0hZJGwbg3USLcVYrXQ28ImODKNvoMrIa7ijQsnafpRM
bSGjhWfnzRF55pT9ziHtYS+eg9TvWaxqNrdEsmpfJx6PGyKeAJqu1o3sAWpgnXG4rkBxzeH8XZkd
ksoP7pknEQj/5yfnsvsVhl+RPwDcksIK6t984RG1DsOjP6Ld7M7zhCp5tTiDrF74z3R2N+IYuFLc
nTWGNSo49yZ5gFEI5akPO2s5/RT/AwSspIyjd+naGY4yUGCKXk6otBAVp9XWJ7q2XhTzHZaGf80r
IpeNgA5P9uO2iRHaiag3tTTiIDVIdGISwa7YMGAawXuVG/zLx1BVcgFZwGbVZ59YBDm32SkHbAfl
Rut2Qw7hG6l5ywgNcuvZoxVL9DPLYFiMlJtFXX8IRkVMaMVZQu7SDg70yj0kqgbtfgkDn5TJGUL8
ANBduPenPdSV+KRXEV2/lUGSDf4kvLQguhGcpORydIrNZ/m6aXSY0Yk4BeZt42XUkvmhhRPoi6FZ
BclLbDK1DqjxI8ErL+M9z3Gc7JFn6oe1ap8LERZ+9mufKs9cwoPa8oumZBXDlhJskICNcRCmVLUm
8Td2P2F9mwMUwzZ/3ZAVpI43abCWsGlP/lLufHLg7p40gH93r0gg0RvUW8E9JzaFTyT2YRdCM9Cr
l25dc6ZN9FYOjCMBKgrTETPBjhAeX8sUEwMKaBAeENhxmB4+5cqEXLuO2yZtEUvIYqGlfyLD6k+b
SB/lZt2BdpIT+N41ZiOHyVuMkLA2r+HzJ6fppcuGpnedKMEpXRMzuVcEJTFHmFF8dmpzvh8r2ejC
6La+e1AYOjB44MCu/jzbziZezgR5tmbGkWShpUvw+qppPnuWITeHGkfrZPGSugqyEG5uwwq4uuai
Ip0d/jrFted7ZA1+wwvhjXvQ3s11amOaYuisGoDquuYFzrETCZpEE3XBhEVC0eabrC+7B1UscBOC
mEGhup3TDfgIQta7luf7/c6/9F4SSqh3c6OnxnGZtrPFqU5c9f6EpQQ2XMfwdTh7ttRmiAQHB15A
Wu2UeAhPEGnoCDzWsmk0HZRc5FNiktqs1RYorXnCbrbuFpGf+yYEjozUMonRl+N5/g+QPx8oDAqa
8RlRAZ7wARy9FOASKHWgv2glqApGtGK63zrL8kszZf+a7MJyvfEXkdvn+xCrEkyBp2N5j8mGDvka
JYJftStgERM82GX+cS6+zXumkrSUaDBtjdYDa9aBtT+tAG0x9r1tKBnAWWqSnRFwharYv7CSQEmU
wXjO87wqIC3n5yRuyCmSkCsWgUtJz9SIRPCULasLyD2Xji+xOkDD4zXQwsvOMG19ZUTPhhVKSYnu
Z9TFhXPt31C1x8YddKegnfOowXBEmC+hrKuKIxTlp8JKHdDaTGKA8FoNoPjI3sVniZ5UJj4yctke
ewMv9NTPibrYv9jc20ViOdG6FyvLuo9tGQtBms56fvHx0g95lb2QL76QHY5XvPTlOr8LNYsXQxo+
xnwpI7n43nl1OebcumJw3tubKUSpuKJArOR+W1mCSyigtI/NuT7wreUQGi+6uzxtCWDQSAXNVd7i
dSjJS1Z+Op+CGVa8x9iXxOXYk9ve/BUAymqRv96urGFPW7bClQZ8q2iEFXLVKaGgpP5RsbDro7Kp
WTakJpAjawlBNuTmriNtLUNwD1gpXwUdhCWeH4+ZOqMXPBAaGFkzRNjEmWubx6FOPBKv8j0WdZjy
NzOa0psR25zvc8UWRTrBQh++k3scPRXBv73b7q6VvR4EZqTu1rNvzLj8wTZGbTiuFHmHngI7jHfu
FUm9Plw3WVcwDfUFvvIExi3np4fOnSzPFNzX1VSkFM9Uv9/FyIDGRQW5EhWbXQOeFP5Tb1+AKOIv
JRmtw3j0ZpDwPsXWW2HdC7OdKav5Rx/2rB9bCq+gk2a3t3GhRZjnmKtNZAN9shhBbLbP4MK5y52U
u6Mi7QFS2D5lTcnARm3FAmRHP04zTZeQQmGZ+FZq2z+mwhpKGLJt2UYo/6vSAo/RQri25Aqm/OU/
Y6XXPT1DP+bnaL/8+WBBhXEbe01gUvomtgTeuHmYlnR4LLpbamZONEHGWR+PUoVlgnemlvuVaI/g
6navQRIAhwCWq8Jdcz1QthAefGsDQZcm0TUR3QHa9Lg6MYJ3XtHJQUCQbtLa56rfdbQv9kajxRBH
LjCgByOf8E1YhX0XyduJqBOqCX3IhRgpy8Iv+CBnM2lKFTkYzKdWT3K+KTPVlPsdGIZ7By2tDI9O
pgUHY6r1RAFRwMU5ghMFXftBSiyohF3uMU8Uxtw8s5tfGC+4Y4YGjY3OsFySzBs+IWETK+B9+AYB
SFd4FsACtQK3+hMjG6UK+Zf4tJq8E8wKja22otsJA0ArxCliEfDT//NOmaoeGsGMqNdU5obzAwM3
bAQZZMClfy/4IFWgkvrdrfEz9iQAXU2yd376osRv+hG7CTvwCz3uteHvL19XMJXBgincCG7FgwOm
hGdTolx+TzsVJcOQTD6WnEza/9Alf8M/p1eFJV2Sbj/ODZO7V8iIibazQ2vvH9wB0b1Dx4gdRtmv
uz85m9ukfumh+iFBrcUTYwgGDqm/fECrak/mOEBRNnZcaoHOX+XoJcSdM9x1o7fQhcj7nC/MeXaC
aKaLqFrFJqdIL3Zy8mNPoSmutfQNYge9x4Ib6MWsB/KO+21c1L/wPnVyoyQVQGGRAhL0eZEBfTOI
WYsx5o3iUe1Ew8glOJDug33RlNDcfN9x06eKcasmQVk1XDK01aPmY3KooJGnkPUMXCUhHcBcEhxz
yw1OFvqjalfEZtKDm2u9qC+DLj67HIMbFPIXUdF5KLOL028OvBtP0KHeKDesUdA5PWfy0rSm2qHA
gS0eHsavFypVxuDZ7jRDKxvxwRXZmfKqcXrGEffViR3A8hGTQ0UYCenGDUphl2HNqyf8JRof1HfN
irjJlziQuYSjL6HCfMHNKpQ20UCqkmrKL2BqlZ4pkZITBEyTfgS3IWg5dURwlTC1Anw3JyGFjKzp
T72JI3dApATsFHlzjWTqW6OkE3UVH0/Fsph2TouvrRSvuNgzIDKrSr7VA46ByqwPnLx5eqepN8Jj
ECcsrxv+9/xKEhAycsz8U7aFKky7RdUUz0vRrvMjB6tqYO/xEapKTk2PzxV5Gje3/4ocWOA0FZr5
Y3dcmyxIfoKjA2mE9HIUulUM2U5F1cD6CJonXGOCVVnXsV6+zmOUY3O6RElls+S80gBfiLowNgoH
IXBnYboVBBKckMk7fxyBmeSdWDgvrtq/gTyzbCtmnsXMQemHwNrKtJVTE31HkmYI5o4NfO0gbJ5W
ZNUijixDLwo0EhZ2UsRQpLLeUEMT0k6vA0wgxC+X4NbCxFVe8aRHToILqiaCdJpn31/TGzmHSkNr
C7C/+i+BBRiuxYoAL8zrKywsceZpTvACiYByuTyE5M6f7nkgqcm3oRHTfqeoQXO6E2ufh8e6TMn4
VAn3lj96dMKKYijdvWyPQvzC0MBU3X+9q0XgJNd3t2vb4Ua2XCNDESq3UoPf7p55QO5TbMlyz+0s
is7HeCV3RU5T9cNFbmgw8Ilz6RZd71C1zADpU9j4IM9YwzFc4Fg+W29ZxqY0w1MCUyu8Prj4Ht9S
hSqYbWCI1gE5DgnjlzRwKbWVcsoEq+k1jZUVfMiFw/CTCxHsAJtZXRZqB8tyX1bQdq26wh8DCgAc
PGhiWsdlG3lK5j3/FdFu5gNqoKEB69yvosfbjimm4o6eEOYQmgH+gYraJ1DuQuqReakVy255fl48
cSOPLgW+Af58CxIkmaeFDfbYP9EF7HDtp59dCTxB1t1TwLFqRTx8Hf35sGFIhnUFdiPpn9Mvvk9n
sx8gBX5S4LMNVTGEkMtu433drs9caK1tGHq0rq7ikRsxXEys50whxRyPACxmWNZaTrmfnZOmqGxx
aGSaQIPW/yTMS1qyV6FnZukGzyTSPevQOJR02ayHvNCMAYUhFpmxzkITtuCE9aOvESFJZhZohqlq
Zo4vMMITRcW2kIR3TVuA1zvRKKfa7ujf/fh8QWfkWXyb1oxgPMam0E5xGI6UP++KvaiExq1yeZg9
PrM/2IcsUl3JbFPzfrQQag0Ogob+9909Caex5rYow+LMh/mMhC8UJeS6uORgqyj59RiG4IQ770Gs
9vYUqEYsNN4W0qLRsCv/XIWnXD52k89zYmmtdDFFnD9C3B6296BxaulQIg3hioUWJ8nrK6fQ582J
YssyCgR5Jz18/Kqu18qvDnXi/pWdHn+K+ldQhRfMqii1hwO+KXWPIApkOLo5Rl37EaIyLwTdIsDs
jFyg+WXXRvRkhUE+tBI8/BTAafmgP4Ljyxcf+vSlWdw6+BL47G5qA80D1Vz4mDnyZTwI5QyifFAE
xXcyb6QrQm+kGpWDyJORz6U0RoHwA3jHZd/IESI6MEo7y3X7W1xF44yQHd0BdOBwkGAgMaqASeux
HjjRRhYJWAGgMUHHETgFHs1FW5yw8WGlvtL4spoUpJQJP1t2qduQ1JZhLr1W8Bod89rtK3gYxsiA
Ju6fySRC2ztDHU0DVHsNW+5s4BqoZHrIAGwvdgx0NP9+vCPrH2PGh/O683WBP5rbxo06UDC8g/0a
QSwh1H90x1pQr8Y4PUE+LebUW5GMaKmckX3MMAEOU+oZLCeCfDCJG6rXELZwXlfqAtH9vLQUxgKY
dpZrWiPrw0IslHraJP96ZUxgwrbWqdcPox2JEwRejsLFKbuB5GuKcoy8dZVuoFethdLkeal26ONy
CHGhcKqzwL4A6KXTCs1m18/F0LYdxFGNwsX/ZTV4pe49fVjTZEwvNQYsyw+5iCnxB042b/pHLnJa
xsFnE3ucmNcIrz4RyTNpoNorYzWArA0ROdViuvs7mZSJdpWQIn2mC+uZ3gqqXK21F4dhyM2ZHa0M
s21zS7ArzN9j/5JO78eGzaweZBFvTUll+kyXMOGJKAFIIm43DLP2KK7EyFmGunQt631iWcLlOPr3
mQ+AYHqD6hNep9k3v1bvjieAd6qnXriW+4Y0GsLz9qv/tjjFZq9+MlF/ZEdiXdmU8iHwBS72mKsH
uDU+TeIAiry7E3GqXLN9g5wozcFMQM4wuQMvCp43SNmDFFKsnZTPrz/t86GRdcHFexT15hZZiwSx
kEL6YD6c+eXJKzu5KQY1MXYKHfsXp0W36VKbaf03fs9BR6X/i92RAZhdFILSJokHh3DgtG1ImfhE
re56Hez1PYIlvmX5Uk1zZI6DcIarS09zHViP3lWso/ug3GRLrBsrYeQ/oNASJUMoGHOfNmH7lwR9
S1ybVi3YYPXpHIJGLWUKky2z06iWAnxiP2Zu7wYzR+OsMQjsPk2jXfRKkBh2qbV1xi72hWlPU3AU
OrvKMEI03FJuyBk2MZafeYEYd9hukLgrhbkoEgsqtfBPNDy/7o+0XW6DwT7K1xJpZKlKANhTeAHC
ONfvDBiIALnPmchGELZ0U3o/fO2Labmhu8ol6Rj4EdFcCsIEPJBqKfymoYim0OKoPALYR4nKBFuW
6VkImIqTp2GlaygFzVEUte9tmsVOx+w+O9mEV2gkGqQCaB6aGcFafqYE4ReAeQ5k/U0fnhKK1yw8
1KeWPxHMwYruUezgkH4H4Z4ISYtnZlKGnH1P43ihs0mTaCfovgc+WfJmFOtg2Co7OeeT1cJXZDDY
92EJrFE/xbeCgWKxiFQR0OhwNWhTf4K+ijuS7beaZ6rzEQGPL8kWT3bckVp1gCs3Ag9KQPC2XOTn
il3wtuXtYleg7Zi+kNe1RsTjxU2jm0D9xS4ujFe4jijT7i+2z6lZFdX3/ykshqVbqMtfmlSbYyno
AaOBKgC3pmDPGwagr0bFKo2dyU+XXMyY+WS2zIrEODwFfE2ghZm1eVPw6eHR1kriMcSjpr16fkVj
cH7GUZBtWxC82Zguw+zZ4h+1UaJLCmVt1PSu1NJFElSAa5EsGPHvtVWRRG26hqi8xA+MDwfimOh0
ptPabC7M63s3t3b/k7I4q62m/4O0jgWDWX/2MuynJczfZ1ddprhMB6fLEsHWH6giISBnh80afXyV
EXJE9OkQdJdISOquMbfJ0tOKt/oZXwjDtADLvkJFTkRX/JRZ53Uj5450FDaLN+qi8bYenaLS3bHN
/Gq3j5ZsUOC7T4ZkhkCjtTcou4lJbkRFB4jYR45lu+4RXEWKsGoV2GsdIWvSJPGtyK/JGJa/SMLy
Eu8Pc2Pv5RP/tf/ieSQv8rKNj+OD8rj9XPVuQ0JJiDgfKnTTjLNTtZ1G3MsmgqyYZGrXRLRuPL8g
x4Kx8CTw9sjw3GnPdviUQ7ViutDw9KaJ4ctL/34qVDcEjhc7HkO4nJ3ujXJIPSrVXjPIE/fnrGi2
ul99Y93w8iRGRIJymFfqvKp+BLO7wuqr2ZzrGGPQSRel1darNj1LzKMTD3k11BdjrROqx9OTexwn
29jS8QaZZQSRasTADW7XyWYXpywni+1Y7F9hrkwqGaHcXUCz2oqtA5q9/54rrbr5nsuYYFvhscmE
PaSOfScNy2ELlullU4BCpho76LAvzHrdpU1TIjLEe2WaCZgb/fyFpW0utiiSy13KxX2BXTficqRS
qkij3N4RMiD7HwlMMbjJEGOl3sLBqi/ipboI/MjRnygts9GlJ3Lk49tfAq/dqCwpJ3B7oD/ODeN+
ZFd7ClMEY2AF+4VYy9g0JQvYbQtxucgOK/iNGK2HsvS5m3ew5vcwSSXdU2NbT83D4CTSOh0o0uuO
bdx4BY8amiyRxBdbsjjC3etP/cxXS0knWayfgRzg22wb9hVMFmDkFy9xfBF3P1MF3sVFLVZ4bBJh
zbVtrt7LN6d1OFy0GFC0093d2tTR6puw0XL2jYXYRs3d7J7035LZgFHpmLAqL1XIngiSZjBU4KGj
FBmxHHKSI7YT0AyfwGiSOuplLhKqv2NxEzuhvRF4fFxEFwnK35Hfx4e7LcnGFqo/Tf79GcIzsZt2
IkbiMF9lIy/400hyA3fFfu8yCR4n3wIOsWlr8JkN7b7z9lgZhG0ISHOpCzbYmYB5hKwCuFY9dNAw
eT/4As2CdzbMB1at9lF3Dh6mjaUAkVY/+rTL/Ml/R8bfYi6Hutfw3bvXgaXa2t9jts+0JY3GPKFY
qt3yM14Qorzgh8zoSIbY3gSjx9SJfj7CKyCOq+XgutpRs9exe8EJ931MRogXm9HNDprgLBGlUvSD
buHFg8dbfn31R104RaFjWO1kfVwYeliIIL55FYS5UcrZ4uR6N6W6vQaMEaPTUIrV8bx9qcPdHjYg
gSHupZEBKb62fRo/Iy3it7egeF0OO7KlUCkKwSVlUaybi22UnZa6c/edHhDv/WhWpjdqf3DYd7Wp
6u5S2u7Js1r8QqmpC6svywtrPHalsb8l+wbkjNtjzeQ+IaslDx7wvOrBCw0b2F8R8SyIbsoU3tIt
jkcw97g4a8XWk3oFzJ4z0z/ZbswdeGvAVYmsmyvMPnBVmZ3J5LFYZlGZ0q/FECbea8w+nRXyKCAW
cPMmTnu4zmfVOa+Ykv8sR1db/DdZGCNg0nIFm/Dhs3AbosHp6ugzozbg2ftyigq/rDu/gNJYzLX5
yPsjPJ0ZOKYKbRmbBdYh8BJxYtDJkq9UVUYaRuUnJCr6l1TVF0jiVpdNpzIQYQDBj38nesLtIcIB
XrOrhZGPvIC6joKYe1t9ttelFlfbO4qd1zpQNiqbvcTsKj9Ky9VSROcfKbpInU+IYEIZ3nrFruJo
Lo9hqWeFzHoKWvzOi22Ir/eyMG+2C2JGkX++hIUJAIIhL+nOAf/bVcK5il5D5eoO9ICtn5w+ebMh
lij7MjO/QBDswJEnSC4lOytjw8wkY7TvVo3+dIGFZpJo5HMqQKybLGKlaP+eXIAHzSti1dppxvdy
ynR5sZfijzDmYGnUzu/VlDo6OtVB8DquQMQk22+NX/4tkLuNQised5s+TAyRXlGcWBQPEsnKXylW
7vqC0Lr6GjD5LE1RiIiNrsPn3ZGhJkXu5hyvfMdA1VFk+iwC1D5En33sOY5YjXlFxNtZABiI/YzS
hMQ2DPqRhQ+O4Zl8hJLiU17LABS1D3fUSKuA/IiaqvAcmpuiqj71ayXzaTCz1wD+H8aX5m0gML0u
xzk+E+vrLhkp8rBnopoFEqUjv5wcqTHBksz6kX012in47TntK89zGAzJxKJU94qKglBsaNF4b7R6
nYwCmkK/yhpZ3yzVVQt13aypNYBRqA5u4iCPAXL6UDxgiRK2snmYLmK5PhcTGgfdHdNmJYKpZpNT
L6q/Z2Ja+5ZVk3qoqUS6gspjEBNgMKyYARIzG5eKL5wqAsbaRA4U5OPp3DjdaVB8HLnHmP4Iuwis
41913D+yCwXaTn2OzCxe2aNA0A0dx+MD1sXyAut+kkCIRknm6U92z9nDTIYLyy9cK453IgApqvzK
9RqVrFtmpquTMoQvNdM1tFNV0+WoIIuNgBPOzSgYSXaIkD3a7Xagf2IGhiDACREOyDt8spMNLtDn
nTHeG3z+0x71Qje268MNQwMkB2ygiCmwXXQiAPoIndq270GPbe5J0s8cxetGKD9yPLn7f27i3FsV
8y8J1+ta3X3aaI3Aw/GqyA23F3rQGcW7FvOJqt42754HIZu46MgN4CS+Spzh4S9JKz8fFMzXNiRq
RYYJWuKxhXnUVOq+uko5INtTt+pqs68TeCdkO67G99vSs8ibwYNZxd/4NprCIFQJn67zeJ812iC9
Ss6D51ttA36PxkceX8SMrvbNKOly+CC/jkZiu131kDLiwokzxxhNjE/qQDcYErXIzK1uHCIOz+n0
q9c7+mz3aG0YGdZ1hqYAAVCDMxbXXW/uFVYVNocseQ1CGsc4bTqR75EGqIWFThXqFfUgWgys/1gW
2BjeCdb03/WkqDz7OrBItSCYSQf+CJ7QbsF8pOdkvXKKS3+WsLAbkB3SDsjei4nIrBOX7zg8yAoG
uX5HmByGDpBXF6ycO08Jzpuzss14t+fnV2/Av/mi0bhc7qleYQji87dThofHKP3sk+0yXIWp/u7i
fdNX82nHZ2S749AlTIuR6OobTiflatpGROR7gfDDHlehsJpgSFhzFSaFKd9CKjVPbT6R7p2u2DXC
8onTUtypqGaB0bpfz1G0g++x25wy4E/BATop4QJOUT1XTibzHDjbdOSTvXn8/L/z6165ENBIpUrN
oELN8xHDQN74yy4CIprJvnIq3WXq9YxZ9jcdjsGZ3FVzMdpi7imVQ0BWGJZkNbg3U6i+YYO/cqTl
N7+gcR9lBm21vnl3gpHYpeGgLr7/Hl52jbqiXDLBgxtdtrBhDKBGbbwJeET210QlHKLLNxvsgiXR
T8T7ZvfS6KF0XaNqoMkaBifAn7C9AvXcMD6LKYKx5yN1RjfKz1LAVJw0lDkNw+Nc2EOypX1qV8uu
ehAE/Lz0L5ewX+dV8UtmobhD9RSoeGBus4y/ozD4TS0Dxvo+5iONd/07MJ4bp7cuecHusGLc/xEb
CPlAS0T+7t3cR8U0vfcvkofDXtSbio2cC40aCy8kGhVJ2Dp35OoDH3epYkNMzTKAJKq5i2cw6f+r
Z8M7UkJ+PF2NDnBtVi557b2vQnABQT6Pe4S5UrEq/GCFhkDwhm/ifMdgu5tL/GGp2pT20KceGRBe
7hKolHxfKAJ5gwjlMIZTzANz6amsx/6oakzHrtxXgzIX2ftWww9uQdrlRKjzj3wZk6+xNCUSEuCw
LwqCLs1R8i7mizkF/vbLTtZ1Kft2YaEfr0TuGmI9/I3dm1sd98FOhxi+tA7K+5oy9AC4Ht3HEnUp
7siBHpCVb90ozttQ6vCIaxRVKe9Gib4INGR71J0MIw5dSc1YzXsUTXfMfJ4/YTHD3Z7WkSBkGFAl
GNrX/Q7ogCNWYVl6sL38/ZLT5YyymvlxNmh+89/8tfPMEzXZvZxnNfwIKJ7yxZ8x7rRcDv07ftWP
NBWknEaMpo/LsupR16VCEf8NhtiXxQzAAyt5VXpbFo/jM0sDPUHgqZ59tm73saKKEx+0DbmAkbWi
7dp4pQfQ5JSHT2g0crMlQRZ2JLmrPekVAWtTkItDKTrRtr8Ad6b6pCbJNlR5zKmq0U0fhmqs6Sa6
VAFOBUctUasd0nBe09rtNJ15d0KQzSTekcnaerdmpHLeqJa4CzbWHdBmDEjhjheS1oc/KNr78x5a
hzRi0ySrpD0eNCoYK2wMXbVfSe7pitcqOdFvr3EAf0uUOyNeZDgtbP7TYSRunPP+RxaqyKoX3xn9
k9/YmwLqbn7OALzSln8/Zzfq3Biyr65TyUyp1r6xdEULiXtOXOB6URgjby0XDQDFctMlzUU3Oe+F
++lSTKLfNqMCCtfnLXEQdcSlyTu8neBXbUXnXKrvtzpSm30wovJwzoGfmxbhigALBrUA4daYjxl1
A0M8beCYptoHBvbw1Mi9gMPp2Bdi/AFCe1+ZZcu4enYuAq/zyv9SthJbQuIpwkJmQtwQt8uAod4J
+pWajq6PiVW5IJxbS/eaQf79wI0ii7n9idsVLh8FTgfqUb4aP8BLW+G/gij98lSufPgmt8pcZTNq
cKRVKpd0LxeUZBTj3AP0mgw28D2z1OG6Lv9AUPwtZBu3CAP5c6EPbRK65L9T9E4283W3HItb0/7P
hWrtOnRwOHOnJgK+MtGMiWtzv9Qtlcr3VpUPkCFYeIGtgUYnx+ouZKG7FVS5SZ0Ye76GS//Yiow1
ch8bA6C6YSpjk+Ta89pXdxcZUVK6E1LUUBF90PIyw5zI4wnv8sJlYAOpMnLWAbCgRyzFmr9Puu6S
5nUsVpRozdUpKUsjdoaiCpYgVNQxMZjysJLWtuzwMZOc+1Kw8vt/kJibNE53jd99SctgzXXy4REE
5SrbMf+WJ3WCM97QPhXKN1r2O0UvZwyIeVDbQ0DW/XopF2Hhrfh+D1tUtHtvaKPM8Vi1G8EGg2YZ
T7Gn4e95v/diWBhftJs1kegnAsApkd5o9qE+KkR8zoOUcHLc5CXcBvIpDGVrmUpAlQiZJj1TrwRl
tysTuyofBRfSDbJJVNvFgISNJ97iCeL9fh4gRQHu0SQeWtH0UQw/Qp3my2Nzl5uXeP/x956zCJi1
NRfgIGs2DrLaruAkfiddTF+C7FnxWew91U9DEw4CSDO09wIMttIGI2dUA72CCP/OjMyfqgp53NXJ
c7k9dVuPPikszJT8R/NgJHs8itA/Oi/1QPTLl/KWa009lLPe4CLjh3ZrLa+rPG4BiVszdhFDGR3Z
glEjSY1kG41Rio3DbZ4PHQ7gZFh78j/o1Wlt2oaDE5tvF2GE3qMlimkLjNS8efvKClRxTAy7RbhH
zFshCbO0Nxpbb1KrPzeko1izw/5pZfMOWaZ2DMNWKmxOaPQZF6yq2ClkTa9K3NExs4TaO1rUMFwQ
p+tVcJUtSMyogzzbDR/0Zduf6hervTpxWqsuvVDR5XcO/bb9c0HugJ23/BhtkXPTmbIVhFMmv1aN
BlMiaB39FA/LC9zAx0Bc6Pw/i82wwOMMZxPU11O5VYogYO77JAoiULFdoqSzjCgoX/6GHwHkYGWv
lJ9YTuDb8UEh4uGJ4p9B8qNupqhjpyK43Gtuu0QVizB2MRm1qHV1Ot+I1AjyoplC7KdEOLFfsoy7
HSlqpVGOv4gUOCCAWKtWuTsqHMxLLUDZnWz+uM2CPnb1LnVE14XJa7mn4hKBCSd6Uvn8bmRZQ0Fh
2VR7TA0QoAisdchNKziWnkD0yPeWd13Fa3a6qLo3llkgO6Yp0vXY92NopTJUR0PmLhktuHou8tNg
cMeKQrIVCIaQpX+7jDtUOecYtj4H5RxG0ANaEQ/cNoBsK49BsdY6kLT0SM7rRcMRxu5GewyWQ+W3
9g8ts/b8ddUFv2X6g3CVSePW45HOcbivhsFFuA++/kEawgzTrUOMs7J4cYG8XDEFG0gaaq6QgzRl
Hmjmb/WcAUwToJT9u6Hefy82lhGZ7gEYvjVmWGISsVL/zYZSbqY/TP97A7FnvsG9EfyYFh5XYi9f
FHhRslrdRHlLu6L7Jkkt77DT5V/o1aJVaqWt2sHKwkoT6nvGfYHMV3I3soXufHWa3xS5DRZdAll/
R1ECRFqTpgnl8jbLQiL6Q0elwouvkx2Ft2+ablCcmtt4dxfMTg3BsYNlr+LWTWh8NFNJLV1xJWvU
LNsKzS9OyaGXqBGsMNSncVpGVA74YD2xs5GULeWQkqnKRy0YpDYGmLuQUEIrnzCAFdse6IbWL7Qr
U9YiHP45KoTkCyxVnp5h3F6q+ptsT9Z+AP1Nr2Iym0G4w9dqcouVP0Co19ddPP36pjmMnkvos6B0
P3GDpQAJiFH1CD7fmGmVDFnXKof2+dk86/SGK1PJ8Q+WM9YJffVyLefhXu1DDGES7IDy0Pob31pS
4RGdG1X2kD80qcfHQ9yyg/umjsBzCdmryQJ5VVeFakIo+UU24iC8lYttFPCN+0EJJx8FoE3mqSXo
ULAdMlY8UOrSrGq6iKboV1a+xg1LhRmIWDYlYybuQNPuyCI+RJSsL5YKfDrv6ZpKciVC4fB7m8Fm
1FbymKt+Pj0UAj3ckdfJAw/oyNW/i51kUOLSIuNjTMYDQUokT/gKX8a9IACU6QItioBkbj7hKYWW
Hj79lcrGb8iaAyoeOsDx1SxMd/S/IG46bVvMFIqk4q+OLFIUWWLOMMkPvB2c3l9onl7uO83hKi9Z
ugLer5ZJKLOJXSRgmhMsSvu/TJbimvYTYhaRYAzUDib6v8H/lQNwjZpB90mZi/ATA0gvWPzkBrBk
GQqncMxpivdExi1Q0NIPV542p5d/e41Q6Jgz8H8H0ydq5g8aKPnDW62a8L9hZyeqjis27KZBWNsE
w63szQlvZONpAt05KmdvvB7OKSgTaPpFlp5sp+jJqfbKw+Iasbdeesg6+G14KxOg7AtrAO8U+i4K
ems6sl9lzCHYBwliFlE3EU6NlgvwRahuez9ACvzRxBkMOPls+7EDXm+td9G1cbC1NCSg8Ua/jGMu
8qDkfFXnhgSOiodS+oJf8jSli3ZqNeBIJClia5yE3yvQ6suSu/PBLJh0BI+tbAhhi/gOt1KmA097
U0Qj3fJdOJAD9bzvWIGWDJczbPsaD/UiH928HB6RbbozsbCIZDaRgVoJ1BaOLNieylWF85HITVa+
Tj1OqQWh/TMJzU4KjTkGZlTAfdpCxMIgU/t4l1NLtWz0O7zcOceB2TFXtpvUh/35fBziqJjmekao
srx8s1FCeuRSh4mF9ef7GNR8lpd0czSb3bYPFt9TT/okYmviEPmlrVmVRM9OwayXpa69OACcq6QP
wOsLM4k0g8mNx0b7DX1R53U7K7sI5IB2zM9d0QQ6BCSKuz7MRGQNfK3eBJ0N9DQvRwkC32y45N+B
dPb/tXLEBneH0JyZResIZ3d1Feulc9/bG8AJYeaQHj6OrGSwwdYxTuaO1PfuvhyTCb52ZH+57Isj
CkThR6Yc4F0gcCg6dxRuHIE4ZGu2eB1XgZI1ILvxxKr+YTLID02+vrV3mCwxESFUEFdVWtUoSKox
dnj6mz/KS3WR4eETeTw6yf9DGitZhlrSb8YtlkONQ1SXujMiql87f0MOCyp7wmIBb63kKhaNgj8t
cSbnJROaM7TSVgQLL4mxV/gU4n2ajdykbWOV3Psr6i45r0RrBcJ+FjU7Of/jhMLPU/KYjZXMWNfx
0MtMD02OcjmIF/6GihXQV2OK4URL14PY8FgJaz6Ezo88xrhhKZndY8MlMfc9wrUfOPwtXTJCEWAu
QT48Sc8kGCRMqO9vNu+4EqH1ZojeekLae+HUfZGcvJoyEYz0sI/vmJHiqXN/4tpopgDdVySw+zht
YWENrS2q0HHfuW02w7KZ1Ux+/CwzUTxEVFBGBLG+5ZGfNy6bQQ5YKSzjYv40DF6MNhyJF4dB85D1
16Z6slNpQRRexakOMlrTjqJASJPni/9AMHvuRT7jdOc/aParVBBUMLF/4te9F0rkAbpPmRI7eUzF
tjfhs6ndvv59jF4DlnEcCUcD/XDU4p95jxH3fWIqms8PtW5CZ2vhnHTvK6xm7rJPu1fIS8qzkWkG
8PPVBDc7PWpAU2h7Tnp6mSQyImIeUKFw2xYyZkiDzO1JsIxXqCG+3l+y4u8laPl/eyoNfuGqRjJJ
eIdIimQ/y5GH9YKKKNPHns3fR96WTqiwSnkEqH2o7wCoAc5HdKxJdbriGn3vRvsRomGbIx6LDi5X
xeFxOs1sg0eYtleaMvz9OlurBeTTGsTFQw2wqH93A4oF3hud3QL5JFmHT7g7uAk06ifzVNcnTl04
7/P3EqvsUQdiZS4gz+8lRXi+vGLGriu9CVsGJPNseo5ysVqqGjTHQEa6xj30gSfmxad0SZi6M2Tt
NM1My18J/VCncZKoZ+4B4jPeLv/x2EkD36rPyC0tySrLI/8XeASUAlB8Gx9jsQThgpXoFqFOINYv
VH1YS7ME2u0obtLxSdqOfveLIsHAO8cisOzaOB7YCBOb4kcQ8pqmh6N4t5QU6r+tVMFN5RdOIKHe
C2wvL8HQqtgaMMWOIuHmEoh5L2hqSqYRYxTyQIOSEcjEjX9JI93zkM0hNrPl7pR7QfoO91Jx6pgW
JIB7+p/ToFX7Q2bx2OCUsQUkOKS6CHw8FITXGevNcr+Vwjbw+g/R/gUd3SdUR1yAXpCVGy49/vJo
Z9GKcMcqes1dkG54VRbD7Km7it5AgmVgFmoS0OmPmyP6DVndxbfY9i12I+0e/cGadHHv8/fWi9Wo
mUQqCxliFN9asr99aFTm0ZTFMQhLcQaNjL8gzb5E4ci1/G7NFiRxmZ7Bg+594WzhZ/+7JWkR+E/e
F+sCd2w0v4NAKA8p2nXtetjIrnmQq4hIGN++M4UX3Rvn6tZHeM8AM2PoAq4JzMikryXc24UeG6MQ
V81oQGTp95zerGmtiI2cbfR8vT5dd9gAncIB6tDZqpSLZHVi/qm16xgkLhsVwESsu06hQSwFtVeu
6qa4rWx6Tu4bAReyCB/bPgNZj5/OS2+sfQLur4hZ54XV47rWrWffwdzgJoYQPM0Y6/VEzS6sHSl+
krE4wZnv22L3j8aIceQux9QCM2XMNQTfdjzDbofnnnkCneryGQIDxYIVb2lWQuDb70KVXro+7/qi
npjQNnFwcKIhj4wIVRJyiTHAFr2+BMUPectindwyIp2hHhLQdKpEijazDuwRRLZsKbHrsY89s6UB
Lb1OehYXIRvNb+iZiAQtP0r1jk61NaP9CSQ10KB5cr0A9FMsahBxpfvRu1Sp2MMZF4uZ+zRofIYh
iTsGPg7KPUO/fSPenR2kvnTCcDo1jHuBAVo5xFiA5Gy30Mybyhj/sIU0yykKQGlruavShCxjHN5x
1pSflN0BPINYtEPSSQW6J8ZhFnbGZitKvN4rlZRplwxME84xrK9a/K3AIK6tBBS1hADcE19F+Fru
J0lCayqE3hZVylXAU6/OVbDrkCEnb0AZ7wa5zL8irUmE5wkJtw3g5OAPKhSzQXA15FMXvffS+TaQ
uwScIpfyAiNWJoNhoO54v0hGnFoBR+MG7t2EWsb9cf/phk7mDWHVEfjqPDhrKhg1KyAEQ70FB2zV
3dHjKPGKcZvjEgyQS8s3SRjLXObS1v9syocM8xn1Gvl47FUuI5YsoZvXHCz1upXjYDG6bEgUafH2
QUMYR2TClR7SWjslWCmH0xoD7Ki4EDXxItFP3yWrDzqxRqONP55BpXuVUzowMKQGA74wOo2QF9lG
krEl6EqNnDHFZPc3Q32fBa3emP7R4vxYe49lta94hdGzirccIxs8lZFIUi7wCOCsZz8uvrEYzGb2
a8+zn6UoNNRErH29WLij+ndfcA6dkS9RqCFziUzs8m7tS+argllhec5JBxBQ9eOlAzjgQUfypb3T
EAtB8gj7rIaa5Jf64SD51aCtIhf1RojYfgANo6ET+D4IgFBcPPrbn5xSRBPwHjHayUcDu2WaVDeX
cvsWbIzACwgo97EKK0dyEBavy506q8BN1gYW3MF6isH+DksHW9T8xHHJAvIGg5RqldcjTQFa1eb0
UqKRF4sodgOT4F49ztp4ecFatjskhkpppGZqnl84D227jbEUet5X4fLOfp0DVnrUN9qrJ+yrNhfc
mGHgu6qvn5sk0AD2377omI65eGfcDjQsJHM3cS6LHvzR79JMQrMSFxD8TIi1X4sYYnwa16/1eIvE
hdoZSTJOReBcHwe3IJg2X3U0KN0C2se7VajbE7eXVNfNt+bemkqIcoM5Gh19WfxHK1f5Qb4REWYe
FuqbIrR5UkU+p6G8V2/a3ltJ+3YP5tvJXBVH+/DtrheHl3l8CJFxUNU8mnikMnQ/P70aAregUAPb
kVFIRLctl8jx4Hp/rKSqneEu7Z4i4Letrw17Ij3SljgDuvwhQAzkeEB/lmnUuPEZqhAUabrh7GcQ
Slndi7d14WwWAi3AxNdfz6W7/kg4QAL4d0X/cbkdyQxcE60p7ugTqDPpZcyymimXwnjbFvtxikOu
fhKq11ePogLGoRU8vaeM3f5F+nwgLxv7Xd4ujgBVtQvZTwS0se+D9Ueu373DcjT+QQjajJA9694u
I2Pf5kH3JHZto+qSERWyhd7uaRFDwpxTdHtNXtutj04FfiZpdnBLDtc+o+v2qYgUsBmDpMQnk4k7
hq34yOqzTHg2BjqCEkoGz0uY0N4ADHjJPyL3sjwRt7Y8YG0lyRT9uBfHnu9DCqcK7o8zwf0AWmK6
U5WHK3WHR3ggQLMw6g4HZ/coMU0oDmVzol3NlG6vgANqpbtmHSWaLGo7Sdd9Xi2Dt66kP17u4UuP
qDqJdzpHDzBh/QpSOVDXICszDFUE6wf5lzTMeCamWe4M+fLnblETfd69XCGvPISUIHEpW8c+HWet
CpG3/afOb+AXtYHO3OA0tIJCY3Pa2l6lobGjv7C4utxRpvudMUin3PdUo1bpRa5kQH2Pa7jErQUi
UsK6L+ITgz7f10IYDGiobqxicAdi7WEXoGJsugRASDuZl8xyv/oGmlny9tJm1DWCsyPy60opX33v
1h79RYjcgdKtBW1VTz/5lxvFyq6Flu0YwP488efDqFD4mY+u/OklowErXcteTNt6tmZHJ56IqADG
MgsAeg4+BSXgay7CmI+cigTbcRjDcEEk94udJsRsaNhlWcbEEIX8789kY1XhKLWSYAgcwUFyocZz
hr8lvYk0OS8NHXR/S+ZzMY1iVtvDZC2oQXq2FtObVElz9Eu0EemZTNPpSPZaylZ5nTxBafMsinv/
Xy84ZXIUzBQekF5pL9U5YBxxIeMyD4ZalXLhzzlv8mD/k+g96R0nlYwSWn1DRNUY4d2dNdXIO0Zh
6xYOiXTzqB3AYQ/w4IKkf0nKbHdewQlggFyMXIwiRZzHQ9JeAasOy/aO+tdXOojWvhL0bvJ0M+c0
dZvejaYSIt24yIX5jzy8UARpsKlmFyNUQxgWtZUi2yn0roFWhN6MLjOSo2As4d0NzHs87GWPAJ0x
c23nkiTVDVZlBAVHTOSxCjd96jqSZFqu/tdAq54KG8/ogeinHjCdXE6an3YwRgiQLOYB+YlEJbww
fKe3i/4UH8jjbON7kWetT1vWwVdI0JgaoYsgYa+eC7qH32r2FvW99HrJ4rrXff6gSYsFxIokp6nh
wNOU/VH6keNqvPOE4L5dkQcXjtH1+szoq6gNqoVdkMngU4POtLKbwAP7TUsjJt4etv4UlOc8eWiH
UTbbameHAgjExLSuh2wb1FHwRhD4lKLSSBorBKQ7N/hROVJEfiOFW9pdsj4EBcZMRfeowS2aowcp
B3tPtHFJ1FO+ogb7mc78imWET9cwYqz6xbBt9lDt0wFtCwtUroWbQ6hhXRS1CYIaMJIZlpHKNbA4
aZhcbRypF2zSK2nGmQil/KegiIb5dqhxiN3M0ObsXnzmSBZiF/SK0DI+sTcvIxdC5qX/PEh4cm4e
8XjhUtuHdd9PgU6Rmx7YunPDTl/ueYmuiroGvgfAEcLE6kAVhK/bJ3595SXWW1po9IXlRf6Zry6y
NgqZUjC1Kk5R5hvq10WlZ4a5ALFEEB/iLcak8/KXPr1qjZsz+m01FPFZxc0Y6qIFb/MT0hKFtpJ5
MHbIjQD3Pxjh/vE286VB+qSWv/rNAShnixvrUdxKTlTlxibxv93PNfmCVX59j2u1p53SIZZpKD3y
XgZ/SPNXRuoMnWUShfn07HAiI8k2ZnVAy0brJNTmla0ai2ZpfurfmkG9fjB6ys+L0xg6/+ECNlWb
5uzC6TSOWTl/wDSwkIwCJtiZXynpSMqaecY/b1eSP1QbIuruQ+nR3OYt3Z2T8x0ugvPiv6H7sEfW
EIFP1Cb0FUTCU0Dg9oLyT8LDLvSeS1uVEDHl0xaKM/eqNkhd7xOpUIgItOh6ELzslum7cf/C1BAv
yV1fQxH4u1RMxBcNOZoHUZThmfjgQXeR41VZ/48g4jBcNPyGyJg4k0b4M4KGoTgeRf0n/3Qe7AmQ
uQ/px3zwYrv0sLL+0BZQUJI6YzKI2B6s3P3Gc5PB/7hb7u6I27bcjFXv+FLHrqeWEihP3nqXcz+u
B+Gs4vu/y8E8Z6RBAzmcOoF8qb4+RSJqSOBRLwnxfM8tMzz5K4k3rFGTvEe2YyFcJbEBTpxAZYkU
0LOu9mqOi2fnFJX4g0SbVRTPl4ir8zxFInvbWenKp+MNCvCwN3ad54hvmAB3o4ul6OkOTruShf7D
UxOG/kICZldEXk52ozHVbpCtNKsc7zDfsDCgR5rZAMSbqOkS9lkqIfcvoTEdmW45oh5yzo6DuCJs
c5AcxFn6qQ77RJOVNbrYfIXv3Pl6fBsrsoSX1R+pEJJFjcts5DbgtFsrqdnARvqSqav+N8E5wvTX
Q/8WlQT8j2AKy0n+HekcFIvhqnqzy9FtIY0c6qWvZ6k3Izb/jzIkQqhmgwXFC4XLjlxeW+g4XJ7T
Vae0uWtrOaGj8RmsV8sz6cxFDnubB8OfUFcCQAolJIGPO/7LlStrzIXGU8vVXoyHiuhRCyD7pMGo
/92zmm/0uMJVQ5/9OR15LINcC5TVbN48C60sXj0z7Dwhij6vbLJ9oFaIYdyiFY8YWdz89SioHgRp
EvQF0Fg1anvTHnEf6/Yoyi9jbD2UwFsZY68gs5QozgttrVLtDq4prkBNI1/g+x5ACPLNM0Y3Uyyk
m+dNPvERUwqA9RXhLyj+/y3CWHfNXrfnbsSHA5K1WfsP6WlR2lqCBYzTwv2sW3dtnTw3H8gwe74Y
UBTMOttAX9B4EKiDBcRZWty8Php3yTrn+R4wzIs7dy4Xex7NO6jx1X8Gtk8vx3WxpQHhNOMqsdyY
KqbbiowFk9hVX+AMSlShI6durLMUMSYdbSd58TRzpuo07GlxpU+PNuM4Or71MihgB1wJMfUPnI5Q
xCuWeHtcRPrYk0yFxDnFvGbPxEVhgHCIFz+1x70gKrVWkgn58YB+M7aDh0it1KaeemhpcIwG2apP
abnycpXHGdu/6z5Fyc+i41kF58fAoATuAPrIIlGg/0QndK2rT9CZluZrmOSusmX8z+MTiOAdRicf
K8r+gdY6u673gsgQnOs8sQEgVQXGtNBj7g6gGxu/+Yqs+mZ9fRmgp5TdZS1dZz0dqOK8ApVLOK1a
cRdqyULQk6MSmNrgYzBrlPj81KsZ0S4GkWv0Cus+BlhpQ35ysTblXVEOVh1Afi/QAa5YgTFWafAI
jloWoW6fh/FS7i98NAnOjp/ZODBsX7As2alMyHcPRczGGKcrSBk8ehuU2VvDFoZUsNHk9FBdL5LR
Ncn1Acwyxm+50JHKnRSS27spjvBDZUR6gVvSFqVrGlM2nhvi4TDglcX+bUpgUbLUFjPXBkuquTii
OYAWXYD5GrGg6GMFAuan9A25hLKU+R7ozYhs4c5NkB9CaT73pIDlp7cXg9coYjZd9N8MlAAa2jYR
YFJOeaQjsifcMkpSruKC4/93HRKVp84v4IpPqcJ8y6pRWdobQHESIWgq7vrQk0N/jYyMfAKlzJP2
xXpMWHeiyFIKMyF8it9w6g6gqu0kz5FxeZ33L8LG9F8hzvzAU5dECprk7feVSY1uhH00QJwknFPO
Ul2ge76wrAcD4mUSX1BmwWZHHZBgL7o9G+7TANyYijxrzyDFhxm6GQfp6UUax9kvCv752rw/BDwg
OruKafxPYFwDHrfDgNCumhLLbJeKrcpWz2Jaulswc7eanEjdns9/g1KPbg7GlxKD8I0puGBDGkcv
+oDZQv9ax8pHqVFAESTD2lRhSyXW6fPMGugm1SfMMkjfBnTQ+qFldVai6BTMLrASrEw5uaipiYv8
/6APRx8hQqB1P6vE99uG8q5deU0yIaPSHj7Kj2jFQCkJELbgshQIUhxA7GIjuxV9QyYquwiApW3w
WYo60I84FGlWPUyaGXxRSwBz2PcFtTArGycHgbKt6H3f6nMPRwOK5U+XGhkgZhbvxJLxMCXy2O14
r1n/3avDnq3zjSCV0aY0rwexCbdd61oRGOTYt7xPPMKFwZ5+yJZABJMtqvMrfYLRVAmD1ziPDUHl
K7cbXQ+8y6CVNkJ6lVwh+nFpbPbghnqcZayzbkt52kFRHSalSLqL3uEXEzOaTMlvde8THtEiH69D
VnzdiUlLL5YbcOJQ2XSodiUpZow1KiO+62A1k99cO/cpCaFXS8o2ttEK4eVZyaB1AfHB+N410egC
xMsD4UB/es6/JkQXNjNJmEb0Gs9KnUHxBEgwXtHCSsr2NyrfiUD9zN/dBV8o/n1zZ8PfseIu2Qna
wmiSfyke80u5sA6PukJ2ToRgsbIpk1U0pI4p20fJBPKLao2NU0MyiaBf8gEnA+3WlN6JFPOYoFfV
quyOhTY90RZLeZtDZp8ZKew8bAEr4RvMtqD1x14RQN4XNQiccTcfJZ8jagY4rvv1np88UeUUFd2x
QGTIA9IiBKeLX1IDRfTO3fOoy7qcFp0Ge4QmYcoV0IDgQ+2RmHgelLkGlNz824GSeD51Av3Wwb3+
a4sGwkf7RuOBE7IICirKJFXFN1voirmYb3tW6A7mlnr1VwJStE82jbjy4jMkHJW4VpaeOMSs95/6
lXUIrZ30c+PR/QGSvW3Kba5pdP1tBRISnopOutlBVbjbQiZgmD29lAPbDFhthqWzCdxVdJEJL+mE
1kHTxUbvWctFwG0O2RSJK95pzpHMoQ5kzd6xfw1a7CsULmD9PI76RcCxo1AWaZE/64Kt/pyGlulI
5QHsvPRoIroLZbefDEh1bJ6WQUpx/IYfq8nDP74k+gra4IUrjXJ7hQ82XBLmNBpAzz6O8fDZmb9L
qCepE52t1Av538iQS8bts8gBX7sScoIVIihyx0SXFHJdhJNagQVxFx+R8LIUWLIhGfwXxtgoLsPi
Ih3wXkwARQEbVdzCIYQ4mAE5kwU73Dg67sTPjp48k43dXBDfEVO1W1+YPl+WLcvvUPnE+1We/dLu
WIj7L2zPDspoUwFVivknYlwoJGhRvDaCfJNV0ysdUIUa0opiWpWx6mwfcjyqjmfFh3ZpuPmVy0FG
1D2TucFd79GvsUTCiWLiAHsAOhzoHdrgKeZnwGDml1btlYuia9Db5+ZTteca65/et9BYjyP0Znau
CBeQ2B6LuxzOfIfiaCoq4O/EMpUoV58bzdzTdlJ3UBcV4NvnbNHEvz+KMhi51wqtWvh6hG8/a50X
vr2UOZ4omTTOpvnKQjC/IIb1FeEDwa3xRZSqTBF/1qmmn9pCVo2HA2k/zZ+JC/bCqSU3+LmKS2AB
TfpF9rvdeStruPg+1qF7K1VN6PDyWeLc2oQaFL0P/C8dwv37roAwUIbEyUHbkHJ3rAxE9U83kubC
eFOgR7Rvq3cFTyOcrHs+1M5T7TNrTzgNNqL2PYzJZyCVFjrSYg26/Qy6ULl+h9e9B1BERwznFW+N
KGxUO5MdmdThc3Z33sYZL9wKTqqb6cfHes9spN2dTsiblPusMkHSgnZIeDtgSdUSR5VIQP7CjI54
rxm10O1lp/YgRM+ikCNH6l0lmwAzb1S2Vdh/6ygKYI0QjOt48seiaMfSDpNRdt5eVecKtw/HPT4S
zvJngykZZFOpUUhRDjNEx43Zcs6nbB+1leMRR6wsZV0AXSNoNjAlj+h7WASJgaMXjxMCQfMoZOKT
mIk5P0kcJz0bqdnCryIJII7ltWBwohvIDrE26+rrxEVzO4GKVKRAEyVNnX3JjNvJRssLTroAnVtU
Cs5N3fYTgT69ten5uIaDtxBjCm/nAdDao9lJwwHob2WZ7fMEmv9kSnHUuKfGssJr3fptsUL96tL/
BOXUZa9XCKsU3AKx0sP4R1OnBAUZR69NvWTG/mdWtn8lCSfMa3V2ikrjpEqpD+CNKvZocIL1PD1Q
0IDTPmBFUE/QIPhLg5hLLMjFUOWGKeAXd6lqI6glVXXSwHKAV20WDnjpAjuXSdoeWBHiguk2D/J6
pmsrs0PfKzLv4X9X6OB7valibtSh0VA0dOzz34VlqfQSxwnJY+KOMRpbccIOewo53Qgr8hA6gy4F
QWG6pDa6ZuCMwa3IIvGj4qZJ48SsCmL39UhMuRhAztm6kK6P9xkYdQW8LW4gOn9QqETn1z1jeYg1
IsnW+VACSnbpfbhPVuf1Q+DsF1WfYdq1n8Blgs7Vavq9ZrNU1BG+BcoAUI5kSQ2vw6CoM5my3m2u
MJb/E9Z8j9nRv0o6vbFy/VgAnxAZxXFxixO5rLXOmIQ8nXwSaZlp+hN27oYyEIduWW3/SZzzsPtq
XMAQ2SB/Hy6uj+lreqp8/Ktq7OWERHcJCWANhWsRodIbwHHkYtF8Bs5c/dVjo3vzq8Ka5FIu3qSH
PLLQoPNVBZw5G8N3a/7IyJ/Bp6jUm0bNoAdzIed/LPkHhMgbzTZfJjxgcFc+LS6Zml6YJtCBF0IR
QDVJm4YtxAiVgWAZb6c08vubOX23lWOpBu8qV94uAhitVeEZwAFkm6fEqkR8Ma+r2csh+YbHeEib
FoKwxftdTk2cGAyzNKFqqezKDMjXoaOH66M55vYzJ1SCLYEEKFrtryrOHL2CZhLHrumbGAu3EWCk
ZxpAr73L4/owasloK28wBHmWXyFWa+hri4CtF+2RbIfzBJxzNNys2wDTpKJrUMChcQWEW8XssTK/
UM6IKCVUor/iewSeASeAA6jd8tgC2DcKFiW+b6DgABXeVeehqQtRwE/LcCUBeIyDmwbwL4dWcmOQ
eFzWKlzXd/EQFnOcsXPKOVCNyVXrf1nnVumZPLHHfYb1zs06/JdSxptr7G+lntM7irp9utHHw6jJ
fZTSuPRZECZ5bz4VaX+xwftP3RAD9DXngoHsUS0zA/9uOGHCuk6QTg2nurvhwUNwtzrcoI/oBJKa
yXzCnBXHwD2l9qtMwZtSknjJm6DVoh5CQu6Xo95f20+qte9mz/zgt3NCfJYVN6L9d6zwZsysleCi
2okFGs2LpMcZlC1mmXjNAzw1at3tWNT391XYlhUowZK9RSon9xEihg3INSYBgNKjSeK5I4BtgdHo
KvdV7qksIuSXQFZE/OKWRWbEQk7TMlSQpNhsy2vXw3a3HZuXIJMz4it2rKtsFRbIpJ4uid5WEbWB
JAkVwCb8fiFPotVeD7ZVJFxp5vP0sXfT/d+UpiTAxDvIML2sThdezDc8cm8IOY7qkoxu2gIejiw7
zJvtVsmiKZBygfpwyCm/rVu90UM45ZqNDmpj0Hh6KPt1KF8DzOJDuflu5UKRfUuKciwMbFi2Y0k6
W9/S+VL9KE+W1Q1DXhwBzxnbugQNlfv+HwZOkD3H3aAnmiXgWKn5cj8NmXrN9L2kSTJjoHm42ukZ
Y1WzfIq2u+2ngXigSRsFxTZwpdJAhCEYT4LfDqEQbc5bmwy4aAqdU2CxiTBCIl8IscbCOrPuKiGC
JUZB7SBMtzDhsCwfu2eO1vQHp3/O2NjBjW331JgzYFjCuAjpAX6dQfjwzYEM4aLq9znQLVzWlPF7
5aNVrvU4TRoQReULx9L81FI3PrQL+zRCqNHxKia0zycLxCFqBhtFluNOHVxZ9n6Aoc6tgPPuCFUL
z79M9VdH6O+F1iplRGTIupWhyuY2YQOk98yAjV69uqn5fIHXQzZAeJ2jNUiYjXEzZDejsxWupAOE
k/P8PBnpvXL9HGX/F0YAMtkWz/zMbAHXRwGJhj2wOWH34I0Xt5lTAyfO0NaSXHwqEayp6KmiXOpQ
aEYilZ0WWgVF3vOEdce9m9Kei9dUB4lrT/6Jd7t2xAvJrQw072IHMgAwbOkATt/SyVQjVOeWsrf0
g5NR/Y1gWDSJmsUsVSsB8VeRtZAQuT8zCjwKq42oC0X1UQRQgpxCg1j4A/bHrgHJ6Ak9GiaQUNim
GNhShsr7bjb7u/wGwYQAPCv0Qkz/cdrnwD6aE/rX+AFOuQeAge/mODst9tXsAbMrALJ5Xn5WRJEJ
1ZFl4DxRLm9ztMbBYxDj9Ad7jcV0Wm8qHO1QbQwn6fgTUO/xT8Ec4PdTCTqNWC9qgWynJqi7+Tx7
sjsheI8JRnIl84OmIAQh6/hpd6rHQxlj5MXz5SOB2tmLr8jrvSW0bGu/eTjHRzwP/miMsu/UgqPg
yu+2aLAElGeBm1Fr75VQMu0pgvpxl8ApWMWmsYXCXmMyQtOQt54Gxwd923cLBXySFysmCuL8gmGx
gdunTY0hjcSIBj34vz2/AzDIfEA93zcXomaxKX1oviLHq61Hd8BA6EBUZtUTu+G2BZJIBBr9paXD
COSjYDYH9YH/1Lty2SZNAjNFsRmEHNxQBCurWS7iDBDD78gBQ63GMkIeR+vKPWBvXjiO5P90CwEm
dZ0X2PD8LWOqQ1KNGWjI8KTWDkhDe23BPHgkWdrttdSCOkqbwqYq6siX1H3vx8M+8L5CO+6+YqDT
l6sfVMoRIWEnGPh/JK2kJvBCjSDkqzgYhkJqT/qWR5vU8EIYlZ3VicL686mOTXFAD4lGrvvY3oJz
0zPi5pAU6iP5whBDvFmGGlplYbeZ8G6/JrVIqoorQh+V6RyQJD5JwOos2lRooNKPg9BOdi/QFgKI
Tb1X6BOHFKHkWJmaRh5sHA1eNE7V4vamD+s4UOwHBD2wtqYiVw0xlqwh16F2jJ9sqOLPG5Xvcn28
bLJm+qpKqR//Zz4n9kVPgo6WPs7aZdKPMQd9ToqX/B5LInIunlq7+9LDgV46ls9xGPVCIHUvb6dx
Eg39t7aEL4fpC3q1GGORROPIo1Sn9iy21srDmiD+VLYZYnl1jm89A+DCE/3OSD9A6ieyfzIvLewx
DQsQeIOE2asIjR7BhIKux8h5lTdoi/0TKXYAUZQ6+0QveCK7A3bl6MjEZmxSvsRuj67CfhqJMjQf
VrZXRv4Jr+5diHpAPfs7/x1a8+2Cg6QH+Khp2UPL+2d7EhMTOgKjti92PqF7io0HpwkFKP4ownfM
Ue4s1SGz333sGxAFGLdRSerp0D7zgecYAVkos83dRKS9HR3lSX5KXUCouVfBMD6qfbJguG0bIPVl
YR8bEKVcA11UFh8An8KCc0I4q2BMq+L6yyC2PgALAK3pzANpD6ugRtYIV7VNsNBB+dgSa/mOhoRR
m6TZr/7NIACIJEOH0jzKGeo7XY6h6BYRc0Cry15VF05ztAHG3FhHs1uWhf4FV7KaBp+i7l5Vxukc
8VDH1GO/RWjTc1irQgJ9dYvp15aHgQlrWLAiiLYZl08+OGVjyMoBeMi1r5s2+Tnomb2xzEEMi63u
r21RX0ZNvCCN8NhUwqB0jzk6YWmM1wdLrgkkjdX4N2AjeDoSi1oscTAOAmMtVtxrmNVqzKpOt6IW
/6fCBZECs/ZNwlRmlm0GqLLzdKbb+1yvFaf+ImZ3NFHuLDaCJT7G9YJ1XxpguBF9mGmysfxHnAQC
2KZWGmisIcXA9OFTPvEhNwzrN8ONWfr2IRor49MzaftvIe1tqhsiI9O1hSQ+nvx2B2OYMZwsGxQV
obLygEFRoCV4xBAM+Xoo1hVwiqw9JRaDSEQZ7ShFFpyVleUlfLYAufVF3QWuTcP84x5Kd9+LMbWZ
nxIFpI6kxDsLGaiDFRR6S6neULLVixCPUK/INuJ/7eqrZ9mRjiyXOP1qAzv6qhOwC9q2R7fOqk+1
jCSeSb3r7/joIn3K1MSjur8tSpEUfSOUNTwxyWsF7bY5ZCPeJ2ALIAsN7HqfIpy4LolIf+YeTZ51
5Y01uIkIMvyW6QLWXsycAZAXvcIOxcK9ZmUjQasyJ2FyF7eRJl/MJFsozK4S4b7z6icW3JVnJSQ9
CGGdK1kzrj4ZnFTusvnIH6BS0gA1jq/kChJXDaBkSsKKf1kY3sZ6y+Fi4YpaQQB0bW5sYQB9r694
OwPAJnJgHhT7gtU63ofz/vEtx7lL+XM9nsxOUhtzhjcDI0meFsyR15zqGIRTsY9cSskRsWhbbppk
BqavgQI9zFjsbYbAZuyAAMuXvzPOspgY8Yyjv+CoYIPMh5KWNo37GAkuFfM2TtyhcEv91HMW6nfg
LqQFzvLrkhmnceOVhhoRIlSqVvweu3OlaPdFksDH57cpiBeXDVVMN8+MewzI8moM+CvUZ5Z7vOct
mXTYcam/mC/tP+licZ0oSvmeWdYZ2m7qDYXsU5iOZUHbF65/G+j4YYm3MHqxeh2fZhYnAQUM9+K6
rRi7t8zB1tVcMWaddST7ePWAwtNtO/V37fMagjs9UQwaNm5eD6G8EugE+quedzUhQPpxOjF03qR/
q3Yr25IWLtwqMr0+RBlmPl6vY4l60+7xFP11tsdGUQhfOwShq+dzpE3tcRxCluOoZzAnoJgoFeaa
tjchFSh1D6XVJ1kdBWmYpTMAVh5T2c7IJMnVQIqjThOA6ItxzbpwwheSxBVUC41IfYtVzAErgPAi
ZV5kE2Tk5ok493siRJTlyefOCGNRoXBAQBsY5NX2cxrN5ghYTX4ePtsjcNjrQnDsYW6qUYRPSRUV
mjpwGb8TwN415RrqAf7SVF01xhXur2lEBRZGCzMVBoduqVIFZtrr/wkliNXR+bfVceEzbHLZEEnh
hVth8P+/BVd8OGyBHSLb2ovBScjoPxXNh+gwqy8tgQy9M+BpIFIqfgqW+ab/4L2es5Z540XPNVHB
SBPEblc85vGziOMNfBs3ay/pfOKbh8HeCwBRV2LC4ufu0Xp/5ifx1xPElnxZD5y+crDsSNHH4TtG
nlIahk+4nCW+sGgr26mL893bHMVEllDeI9LsM5huk+9gtZI3DZ57XwbWXve4AUjbn7w9iujH7H5Q
KSW1b9bcAm8prx9eA6xLEU3qJ68D1JScSzA9YQYNrYJdQmTgL5I8mxgrjJxWG6rlspffpBnrowMp
M6leEIgb7CkYr0xTRJJ68WKrTMdZZECqXcxDtZLUnUqLp5cVkiuDkkJAiZYQIPEwl/ozcO4Yq1xr
N9DSTqaBQ3K/eK77hxjTCeJ63ftUHq06ERizqsOqdj/1rRUQrpXp+LniibgYLPzDx8NHs4DtXWI+
v4pLHfkkq9GCGPezdSpZtItZBSfTigj1RJ9+Xc/+8V801XZK6aGFz3GzCKZoojtugbf6LhpjmdGu
i2vz5RYCHGmq8709eijvyFfDUn2+5lJaheDcoXeebaTMBzszAYVLreGYkVUZAvyWh+bsbSQIl9pp
aow7RlH0EMVarbb78z6HdpbYE50OoKK0tl7XNYyXUUb/Yrew7Df72yyLCM+XZql4gP4xTiy91MwP
LLdIqcjHBZc5sP9FMPE4ipNVNIfaozQT4oQxYnw92PcvPBVhANuxW5Nxe7HuRufdLHgPoQL+ZKdM
bdVvlUdBwAthxlPwkr4qoUSROsjALJ1hOLsm/gts+LcKMDlYxybUOKIbGpu9kb37Q7q2NQ6/SgjV
EkDQb04VfbC7/IVQx1QliX3dcuwb/PY+WgHTVdUukqQR5fpdH7hzYYote9y94FqMJyiH+MmJ082N
x8lOUqzMzdt+prwa25Z9aC7s+DS+v9IrZDZEvVYukVWFV6pjW0kWfijIZ8P1YaHoLfOQWM/iUiOg
OxGgi3jr+eR/I1TrwmaKfbN2ofvqs8d38XQJETU5EqKvK2YwypPVTO+c/7rGHGqlDgX1OafNiEjf
gSAUfP9YYpRHNwV6upGWcaUS3b1g6eTS8WqtT4kJeTzoyGZVFz7U9hri1hT7Wk1Hn9fE9rTq1U2V
JLiGo5H3hOb2Ls2sYtloAh0dC+hmJB1nkcm5u+YiGwxyt2tkOS6sO5svduVqKxNP84Nbuibp5WN0
XeFYCGmcuuF0dmVDffBnOzUTQsi9ktul6P92/65D6rU5p/LdYAdCI3gELK1ciuwsdOyENY7JyVAu
u/2slg3bOkgoMcw2tzojJsE7xTh2snHLy8zQhbfBzrNGFgZfRY4rPRKrx9ewtbCnBwV+stOcbl1N
QPSh5mt7JxLoU30VCb96kH711r+oDdWvEH/ujiEZT9S4UAsqpB2NdNML0n5bZPk557ZRIP71I/BE
ZZ31MMm63VZR9D2n9ZR3kT13myYdrqO44hNOCBg3Zokq0Xc7rW6oslp1/TrfSQIYfV6FAccMEe1P
sEOSDCVLyuPnVE9go7IzKur//Reu1LUm50RR/IhQjHehl9Zcw9Qf2V6V2I1dE1LL2AVlg8Y0VtCs
9KJ2r5HDEBYVESawXAwF7FypvY2NE+hQK1lhTJE+hvAq2barOSWipFubqsPOV35bsm25R6juce67
tD3mem/mEfgOaoU6vd14NmlpzU5b1sxCkGZN5GCb2zyBStyowva9M5IDZv4EqvhxKjmEqnSmh5MZ
rzrZNioAObGvyn0Ra9XBa3UNJPuHQSTZET09HEd7r4pUE2aRZILQvzQynSIc4LJeaJKRCPP/RqIb
wZDEh/rHxTCepaGHy4PDLzQ6la/+catf6U2pFdCbX42AJ2I5RpiPCADFfQAFVwWwTRVMgLXK9X7E
u3SqP+0/hfZ0+ybc018octfyPobZSbISUcTbgYCQ1D22SUlKylbjmYAxk0jRiHBGpYU8T9gF5tGv
7nPbTyqPn8SDIcGZ0trc/APeVyRo/EnnU0KzXxAlhjVdFWYtkRiCIsKZkueFPmhGa7uesqNmEIRb
ClayCrC60ZDOFgB+1ZMv0eVTj2nfpPG3lGK7HgZyDGgcnlUTZaUpzgVAPfoqvFH2weEpOFbEs+u+
Bqjh96RdWbrTLBo1CxMnwE3i426EgIvzJlWNT6/lZMgc9MZfF808+z772P9Koud6ZYJgXgFNoYVF
szDrh2utF9hR/IYZsiCr2be0sZqPz6UlIfBeXmYFerkky26zO4xkCVGCiVArrDRcmgwLj98m6LwD
6gyJPtSG+z0VVk2XNMvO/RieYH7qQmu4hSh4jRVT/9MY+ymeIBDGRl8N1e6LojSaz9CLVc5cf5dy
tDu7u6cZrxO8qSWRWxUCRfLzU+RQJOKabUH2EpAgGK2Vnr4YUm92j2rzp3Y/8CAj5agsiXBa/PPH
LgfuuRMd6uKZBmIGHLPG0wdwi+PTj1FMUX82B+5bFiquyRQid6SYewlOR+aNgkhIzeN+o4fHf8JN
NKXfeZBRlN6B4hq0MGG/KOMNJVSqzwygORwTJDr0iov2qJYio+Cba5h/iychkU7g2Mry1Q+uRlVl
3niNRZXC+KVbHA8DWLjZfHsZhRmFf1M7SNnXmt5EcZWolZP8UnT3wX+70msV8f68NoauO56wa8Nc
/FXUf872R/jS4gm4JYjY0/mGn6PkFT1zAYGzxDDv5bDETj6xxZnSHkl1qOXZb2jbmIzNXCmQ+HjR
B3MTzT8l26O9MUSddjlWqacFHxlut4WtnEHkKU4oU2O3E2uipvcw3EdSqJmxNXC7sdqfRyqZ82SE
4JIWJ12Ynxn9+3n9sXzQ9J9sAoHvBS4WdrJLt1wPPGCpiy1urhCCEfqGKC+OWwuxfz5AEvZ93BpE
3gQIRlIipuOerWIYJDTGbqyD8lJgWcrRuf0QJuAUyBQtDXr5/h2QJ79f0kltYgb8tYk+/0U3IkpK
1h4v8vq3BOV13l/E7vDHvdypaGXDaL+bjJBTRc9egEcPdBgDCBmWhk9SM7xbCykpFqXGQKGb5EhY
FoJj3/n/dNjPmss97RhGh6UR4wo4lifMlDgIHFPwkULa4yohMv0Gs6x8D/U+1izYEDxtfB6W0GzJ
RzUkeoYSAxmw8G8mXwpsi2CyHRfQRVZenvGWs2oqvmftS5m10rJCoAxoRwL5GIXB74ySA/Pcq0i4
qfiKdOyzbK0Lps2KYYHwd01JNdaRSnlYehcMEnoXHDli+up0zOJZD+EuV7NHebgFK6/0BwACzjg/
rjPR29HMPh5iYGv4oAJAYaT0J5bxHpZYR+w6P1b81cVRYURO8fbJFs2YYrMP3NU0JpZUSC6cFbqc
5NtWSIEzma3k5uqlmbKR44KIvofDtK5C2ocMdtz+7/667nmSJQieLLCavCLwBcJiUpVSgl9Djqhi
+Vojkin3yBy12D9zaIO3xdgo7vieajnCPxi9D/3RJjQtCIeaHner2OL44aTnxU00Nqnk52YW180d
W9BKXE3SI0YCLdi3A/cDxmuzrTSNGJtciSRjhJiklLNdxHZ9FLA2+pNTCFstfzZT6eUGBhqpf2Qm
TnzF4lnvrhkG3rFwk2VT2itmwyPkyDfI6137lCZrbNhSEkZye0TsN+IKFuA05fyWgzqfvTOLfc4p
R6oRC7+gWaV56oPnxFc2tHdykp5c5BsFPwXM9+Wa4U1vyaGmIVBGIZ6HMN4xn8ZSRziQoGRmina6
lpLNOvGxs9OT2LL4FRff3sKnW0k06kdTDTowqZkHg4TQsgPyJ53XZ89PI+ZBn53hqH0BMEI+OK5E
tzFRT6ryQPIZ66UfXrkglc9pbFCsHQpYLe2Jp1nTDlzXOw8XwcnM+nIldjQiNaJAVaChguVGiUay
3wvFzXfaChHFtO/hj7gFtZnX61QRNNxh6EciEIDyEZ1+imbL3Mttx0g04Qtvbvu6TflBlFyD4qcK
aKYFUbtsuQb03zufTPzCuF1yDmt3B/mnD29USkyxFAY0a8D6+Rf6zJZkSfzCj6qywVQR4SZhaAGM
xOej5mltU25nlej/00tjf/jNCDMjBPmBcqiWtlSV6D6BJxnKNeKwMPVeu3lBh9bHSDyTOResQiNY
Xi6Hof/v8oQ1ZRT0B1LwEeUldjjnfr89O9/jhSTJ/tsEPRFqxU0g61sc+Ih+Xdd66ZQpyEIs2Hft
agLFdlp8cUWcngzg1IelVmuTZjMaUjxCIE3WrhxNqGo+EMcW21jqrZh3YaHGd/rwgVOuJvq5yg77
9JQzUH1hVVBFnvKmkx95ual6JdrWAI8PE8EnQMDk5l0wB8jHUKGRXdljTiPkBdqZj5Quf8y66Xvr
8P+HBv9iID8faJR48GsA4Ayi6hFevb3V+pTqO2T+rp2aIchG3igpUTo87TA02uu3QXo02ZCjmZdi
obddZUkV/PdwJ427H+Y3n1ziPNuorm7E53YfsGXyRn1QZ1Zcv1cnr4c+efEGxLsd0P+mhY0b2foL
3mH5d1PIVnmvnzQUUam1mD8OWaaWadQjFFv9k7XM8mZwruDC+YREqQDGDQNgtPK3NS8WcKFAQPzY
fvWBrIY/uMGUIAJaTLNPEzJApXKggWAXDxFjqvEXHLh80hAqtjxQ/sq+/9bhs5Dw9q1Lsz4c7xkH
P1i//cXSAGicklpdtGCZkju1+wSJWgwbSlDhAJjh/UpZ+EM8dGoGATrs6GNjG1qP8BRoTtqILjeO
VZ17P8/hsVmAg4MmrhuA9VNMki1ZOLlejm2clB4MODmoFP6O4aovO/PutPOAwUNlf5o50TGQE5sD
E/VNZVc8Pe7NiWPdIjUqF+6oDmOOy3ksg4DJEafDDUcSmx3eNSZeiyplJTgdceQrlrvpeCLUO8Mt
t4lOO3ItmsXlD9ceG3s+TI7Q+TYFas1a/h49ncSZjvJ9qax4t0iCMxEyrsJRqB4OlFmgj5MTuib5
8cupjGHMOVAgMtwNcwOJ7vYHHJwAdFt577pGXr1nR4lQMBUEueqKcaltPXhtbgS8v9//XltyDHKI
w/84ZUL9pSF9Px4huoRj3zdDIvPr8hb+R3C7ZFeqis9PCaEQ5OyFHNl1Z5ao96yfF/dHzCJtDNmv
eY/+9FKAckoRwl8FxNzyFJ8Xt9zAMMfRJPoaPVJ/vVtC7qWf0EJmyPRL7pOMBWmO/69aZZqiAT7U
HpOwyy8B4T9t2fQEwFH3Yn9kDbFHEAFS8F8EegyOe7U/uOR/6bRkGQk+GO+CUbegIU9kIx4GzRH7
i1hFtLwRjW1FWxhXF72W3LsiFPBw542GuNIJisVffOU4CmdJLFGz4Emt2U49EIhOM8AmV7qu880h
rpIaNbNLd9Y9ZUlAtEY61j5+/TsvAipLI6IsGd4mgFqsuU+52jQwM3ksIlKvRxn8Kfaf412HjqmC
0bT1GBCkpc2vb9LwXE6nzI4ZGPdMsMHn1k1Am4OtK6AJlsuKHxxX9U6TIIt1kf3DYubErTm4gO9p
m8RGXPgAzfWnDqIKti7TgySrJbK33FGJOA2YB9d8N6h3OestQy6Kn+BkbDU9qQLaouXKxhMqrDgo
j8esv7/qt7xeIwGh9maU2D98W9exwpMEiHnwCfdkD8pz3dmyCaaYFz80XSde7sX9c/DkC6rqC5z5
ue4Gg06JcuOVLJSENMhG9ORY1nij7te8nbreeblrDNc8q8mjh0gDOeX7Gvt47eiv/Dn20R5Wv8av
MZReQjGFG9zXgK945S2BGHVlELapn1FiIK/aYqkdVHyFtTUpLCCvSV/f6z/Jydx7s2WFeH7mV5d6
1VmjGq1r+zY/j+h/Aspy6CWOb4IdUoQ69txB2WZ4V79WzkwjkVYNzhEpPEdyjMGtTcawgoHCzWtS
lDkUG0MVikKrrcdyqNEAtTeJdWNjLHkAhyrzy/xe38UFruu4T+PNa8ohG27OqAm8L6yvs3nXaxka
XizO7pkKZQPMK8Cc6CGLEC/Hho8VMwBTuhWa7dvFF1+ageo4eN21qCDBECnZvpKdhJHFGiVKHioq
2uj+vf4+miX1i7iZypc4xbRcGYYbS2ZqsIm1O67OsvfFBlmw6NUHr7lg8vgkyEKB23Val2OSLNOZ
wOWSwKg17uMPwfsE8snVGACbwdkSIKazYNHfm40gwVuyh/+2KjU4ECh7Lpnkw6p1ix4uRBz3EMgI
1Nvdpyvtjd27SsX9+8Lu5o7yvazlXl8CTCLQqdRl36uiDzwhjWLa2hfm2tyS+U0Oa74hFGx3NoAA
ft4M86kxRFGd7OK8WTdEZdxs8LpxZ6XtS4dZBPFKNgrU9asXQY5cUCY1mNND2nPuQnjgDrstFuvb
7cFphVdwaJuQg32/46VMZbE3NEjNFGR/EU6ieTZ9ozgBSijbYjdA2jAelPGayRxmtM//eL/dsfdQ
GwxQSLV4UrcSYfngM73RLwO7P9zPJ/GMtCJD88Psg+hpxj7AhGjG0p5ly2hMvE71gE5WxR+B3GOH
GTxk7K4yNDZQOuULUUnQO+SKVPy9++B4WiuUywqwVyatS2kj/xjxHZaJQAsxdS7rWjLFvEpinJ50
SPnShbAeYwZVa9xt8dey+5TmP5ucW6aQ36Z0ZaebPnuXOq2tbOKk1tUgFBnfKGi6O06QG54O8g4D
NTCMYi3+os2Pimq+I79mQeu15OhnnI758/ftF90PtafSgAQqdUrxjSW1sxTsZ78FIoEfg5ThytIW
1WenEipyff3BbJnSJD8MLCeexvEYK5yCAp6ttVI2QBkqESQmidwF/XxjORd9E8Hz3AXMiBK24m2a
erNwrXrxWVmbup+FtzxXspL32g3V88pS280tcQDnRUza6kOIgry3+eTSY3WzOmPeVb5a8q5XoBh/
JgrG8Oppwu6Yt60dGiFdBLZ/XMIMSbF7yXYGZKITL3lW8bAJbjeV/AurLQ0Upo/5Fg6bHU1Rsidb
ljfUguN1VN3JFNT1RSHNTojZCEXsCLlbQbQIMf16UoPEGTbTQJf4rLXEn0F1mZWSrKSjfxHvtqsY
hSF0Om33sZvYCkp+d527zeaQ13z5SVq4vg4KtHc05vRgpxKcmSQV59QSlOOHiCszAw2+fECkUwLw
bgK/gHN1ru8mie5Li6lK91XZs9Fl2VwRvJ4XwD2/yg5PWli/lNiaq2B+nNTspeMzJQ6GLOuPgGs6
7j/7CyYjiCbiDkiWhPyldsaTrz7r/FjnTdHm7AbtdsbkSACVHezGuu7ZGclC6kRZ0EBDto/lYdY9
+Yy4AqKv18Z3AycNRq/E4H9a3u0UNaGBs5yznauVS65Z3GHyihxPYhYzoriI7wiTk+wl9Ws1ZRfm
Xl3YNy2l2mGIujoOQtdpKolgEN8kAEjwCj6JIh3c1Sr0CEhZwSiu6bfu9z7bzCLLummFWQ9y1vYT
gf0aQe3gRk4txlGnVby0mFF/phpaFtp8AwDAf6D8CezmxlnM2TxhWHPfuzOwNSp8xLdF+tAYuKkj
WnGjZDQzYRoj394kfy9v5yxMfI3yvB1QJ79kDtmUe9wO2G7qI9N9GqEPo2t4sNQy1R0ade2y2V4h
B1nE2K1NlAzzlUAY6+2SBIoUTbQWLE2eAsEAUdi/bhcFwXm2dJHYgKlCA7iSWWGLtSW3UiBjXwKm
jAb+VtAzX61QkAFwBkjM8XE11ayAtnr8otgnwfAj2iy00T8kPTUn5H+YKTUkTi6DRR+Xhh++pdZN
R6kfvRGJktf+93kJPJKm3wP33/hWaPkDGOdS1g7Tax6PXeT6qPqRmzb05whLK3n+oSQqqfeVcuHx
LWaJkwYN4xu+rB3+vvA32j77F3Szz+6sMP2CqiFB8t8MSd8JjIlnLEDwDrwpEb0GlVOsTv5kY3T+
iKiGzQkDPBskytyToXHqWHaOa0+JOXeSVfhB7go0DlArVo/HkUJvq4yjSVdoWRYy/FcTdRHwE/HW
S3D19SoY6oCc+uEgL53xZePmGX4pU4/YBCqX2eQDM0IAPvCQms293486YZurDu36XwaVBbT7NqYt
/wVlsAoWJDmxF7+jkqwS1ylwpvIv1PYN/Ob607nYEZM8UWBgVdFvfWywlxz4pzw9Xc/5N9+Yj9Kq
njiIqHMu4AIlbFr9vRsbiEmL9TbOUSytTfkpVVcjh3ILPHxEvau4wIM4zFHXh9wozbdblkOAz4eO
iCw1BuiFKCHNxdmTfxvl0jIsJM5LMjdVVG2UtEPG+XaXvkXunI3mT1mLjNaYtY0hfbs8gwGD6c9C
8P/B+MJ3pvfgL0oo1pQ6FtZ729lcaSTRKH0wZcS1RmLhRFKYBrXBQzIAGMn4+ZAVH1CtaXBXZTI3
vEg+SMP3cLxchSXZdIVRQZYLQOkN7xcWBGbdeTAojlSaqFzhGelokBMFsJPq9HxrOMzw/kG6b5qv
9UFqVR/LEhCLGFDJCVVUC1S5BW0XimCHae5IfAum4ebXOwhpJ+XbFtE06HxdEjjI+w/Daz3Nbtda
QX8J3LMIyZEw2+icpS6+LBijGKIIi1ucsdXjjMWaURw7YiNyxLkvHUk71hdAc8fLeP41AAXR2DrR
thlMRwZDod3fCKiZQYH4rDeEmviZUsNEpNuPUh4PUez2VUqfF3P6aIJ1Fgv+hYc22AWjcjh5Neg0
ASvuOD/wfui/gH2xtmohB5664HwaeIRE0/wBQtAxbjqlfJP24asWJdr13EQNv1+EZTU1SgNmxxYj
EzDrRfjihjCpghl8gHvRroRfiTnG8+f3WXGS1pNn3CoEGRbUaBWc0kvPhv0s9Ke9rpmvXd9YIviA
25/7flP7iDPDJCYGW46xytfewugLU11/3qURRkQQ70W1bkgEHZG9nlTO1fJAB2iojr7vJPD2cwpD
5ALCZ44J/NDKGsYVcIuEL7UviqCGimp4sLTJmVrNwZaNvOYoAiAWNG+Sfv+OSB3xc4C4dzr8AhVq
B1wTegppf+JwOK/j6LxCFECAhhCEwfqyubNaoYA6UwMRpb7lxFK0kDRuCuNZtkuB+byutIQAfbyA
qxWB0UPzVeJOnVZQypJcmIrW0jaVf4LS9R6qSpUaRLIkyThD8ZLdjElWngv/rvESZkK+7hGs89WK
g9s7HwcuQqa1foM0QKWBqep1wVlI5FjwPXCkYlBzt2AaYR8t/YCGfxDa4UWA+GtGAheY4dIcN+Ii
f2sP5354KsOvoAxyqF8YszK4zkDC6k7hfIO0reY/+kjjrdDK9A7PE15MNr0vcnnVagSjfBrNWh4k
FFppM5IZ9MGTIzw5qPS16YtB6GXRiu+3+lZtFmtRcQkwF1+XqeFZ16AeJxNFJGRw6uZiPHXn8JH5
3NLYnqkuwSqWNn72krDfobPZLWfdRywS6rEnFJgeKaQHKJWgkqu3EhKEBt217tshAsut204Vfm5A
VqnR293vSUTiO3C7338CicbvFV1IstyJptrrwRy155FUoXZArclkD1FH9DdtQl/GbAet0ZIXE3RR
1mrnB45m/4Jr5gEqdgWg/RBJJPckZBgG5h64yCyZOAJ3/WgH4+B+5AuHjh6Bybw7JEX/hLatkkRh
o1rqE8iYO+2N/CRrOXQiJB6PM5ClIh8FQKG2CPLgxGcmzz/gMblYQQ5e8pO3mzULxWCz7wqSQaWg
uY0C9gMwCds2fx5Yj497H/QFfgTXr1L/LIk6bfyhbc7F1Cc7ZaCAmIfcklHcbbHT4Ue4TXXWxYD/
9gijafEui/9kho6pZSJNXvag3iWT2llLtD4sM1UaJfXsPnH4+tDPUx4UeINV91GWvzVs4dGfSguw
GmkoWoNRjVMF4aa/4iPEARkUD6JBcbgUnEDTAOyF2lotC+dIzHh5V3DNl4wVkRiVD7MZZq6XJv4R
DhX41m0EjaQaIV6EWVEfe2IyEcoXi6qdnyY+Y7Kciajp2jzbsnqRkX1TLAeRRdbhVNoyR7u4g39w
rZK2SCurS8T9jTyshdxFHKm75X/+qsX3Qh7W3VwL//vDqDAsWIaOkgkWL5DYdqUBP0i5eHpcnLDi
HCkG/ShDwopnxD1s2sdCEAysnauVIwSEHyleWbtD4sGi/NfEourtNGB+k4qTrSikP7Av0JoLdD1j
lfKFxAvQFcJK6oPm08Bf7evQgr7WUEhI54m7IkCzLuzJVA4BLqjttkOMGoyiM26QP/fm4USkYyKa
tlGN0EiEHOetqVpfISKiR4Vj9iRQ53nV98MX36soEqyebxxBOuOtzPZhcYQta5+Pb4WXdstkFz0J
AMt/Zx53fXa9X83BHLcwEF1eyZZZli7zNtIKSir2VTDUlRmfu5OPGF6ZhyRZLvzHXV4vrfW3X+Zb
4Ub8K26l6i2p3OMIY8ixaujhdicmkpL/nYO4m+rwy1KAS/ONNq+N7CHKktplXCIieFoFtwu6y+FW
iwoO1A6lZWsqA2lTGdoeVamGMuIURcnala47wMnaYedzC7kZK0EpizH1J2AKVQsGe7wa+sf+4EiF
YAROq12emzA+7FC4WzCJZ+w5obTY5FNmhHBx4ugh6wzllemVkZI3pRqRsgNpbr8jPlhqyB1ZmNku
fIsnq1cBvyCgle/eqd6naneIT+hzytT+RGantidIrs+Qidx22ryuhJNFTph55Ptj5wgBaGnFs0f1
wfsndPz9+abQR459FXQkimVvOV0RUWPY8NCuJjHAexIe4zpi/FFiWghm+z24yi+Vwpx4qOg4XcRq
qYPVKgmy+Ez0T2Zpf7zgct2pSIM+/r3nYQqkWoUCxONmw/zulaEBTHzh5a8va194OpebOochceTe
znn8VAZl181hMqv4j7DA5KhPF+UzjXs7jwp/5Kq5zyNTRDj5GqQTOjRr0LlLrJRe8QO7I2k1akch
/df8/Wwo33N1opaSNNN2wxa4nEJxURZ1MBtl7eqxODzpMfqhkKk+QvziORJSUNWpoIKSc3GaA67+
Jgf7UqA2nKfCR594unzyevxFyzk/BFiacbbSNbJUIUSbtZvp65YTc4H2Vb3/GAQsl//wdXCR9PGx
v38+A8T2elbFkCQhdEEjHPtj3RIQ+Z1dBtTiqK9JHSXgL4pL49UcVwtFJG/zVJHADCosZEzVdpKk
JC207UWJjf/S43spkyhgOnwPPTBj3c2QASBYl3PDck+LjQ7GIWjNAaFjDCB8XUTdGv+6ik+TZShq
v/ZVXZVr2E1VBeAey/a6SAxpRTiGNhAViyhcs6B/aGWUD2bFlX/mXnhSidwH7nos6lkI7IESHpza
z23njuVFOAKP/xiFuz2/aGx01JI8Lis1UUNMvr+R7nt4nqbjVwBY8b3VHFqjyNi3FGyCDtuv4UMH
hPIorZBG4hzINfkwaeNfEDCpUQhskd8YjKs9YwubUjNfFNuYaYSvh7OrqdWeZuJLLBCulStbL1Ic
OC1SQYsXvI4YKlwJYAGs2F1+qKpEuIaGW+cQrZpZQmcdUEw4tc6udmcipMraTcQgCpoG1L05kniA
oV+4k+s0tAUci0EOuOzaxc8wAWAvisezrK6eGM4SGxzhrYp0wbyOTDjNtgVAYOhM3uolYni8zuSQ
xn58/ls8Kz0u7xvhd3BhUUdxawj2bSNXGcAaG9u6w11k6xAJprwIA7oBOzQjNaRTGKiautzILl4X
CxgVXVmm7aZpwutpbsnxznoWeqb2e9M0Hq9f/Ao3iakJZNyy3r6MClp2WjaDBQgECb1GTPxWsz5n
5i363KN41D5T22nffIN20dRkT1yF7V0gtA6IkAIdZ/Cs2bLbjo8yx5VlWmCZ0oU8c8bzcf/tg4/l
NsPkaUCx3Kt4VmQbUQZkkKCsZXPjMzjF4DUUuOJSI1SoFDtVf/eXaa4XC90W/6oZ0ojs2klyT01/
b2Fc7SUE2XDOrFHfWMUMpzb4Srj4n4VsVHT9dnmtzgqav+22KjytJaNAWD+U1vT4mIJbDAK922lx
rBoNFNFQEJIvqRoLaR5mQuyNw9/MKyZltJ+/uwTLcYfpwf4gI6edIupPEakQTF2uIWJT0uqDMil6
/lunIHlYforwXZRp02KN9S0OzJX+VXNn87bwzndSa3HSNfr72j0vaMQn7B28t6643KQYIMXizazs
6MVQzUzxj0lqQXbd/ew/9N/OPy3tpShtnQp+AVLVRKqIGJj6CFP8dEoDEu1Drg3/pn6V6X2FE8Fn
cjx9TLH11TEXkamGHEHgU8YNqLEy/mOWux9H9A0Qq1o1ePginO9t+oC9p52YABaWY9BJ5k68YWF3
PwN1ST0qkDdaLh5POC1s5fHT8+UqC5e6OrxMP5NvHdiVkA/iFGL7BPi6upscgW4Wc8hRrdzG7CJV
MXvabxzN2b3+UfTRArIlfSSDwPKrs9XtUggPk17cphm6BGn++Fa6jBp6noMwjNaPUjCL3ghx42S2
HMDStJifZWrDi6EMx+JxkL7jEOWMoo2BzI3ptdCPMo69KCiiM3ciIEm5B52fTj3dIjSHlmF0mDcl
HbrA1ph8wdFRh6M8XUqKQmwSs0DgUfZd6Xw2IGiWmjlu5MKSFyoB5nmP2Hzu0fM3dJ6OLcsYwRRM
PJ7VD+/lChJAmSoa9euWzHbLtPOaaJU8zFTSGzhIw8LzVBPmzzIc1Bby+UkC1ABuJ7eB2MQjGQSt
dTFRFt3Jixcw4GRM2Qf8ufZRoYTFKw9N3JSfEV9DPzzAkIgC7QGvNRQRwcR8xRPS7ghyTnDgDYlI
Y++5V6lA6IlN+gw5Sb01R0sSfSdwON7wwnlk07pqm6RmM9N9+OD4gmmFIY679KhY/ZnX3cPV+yLz
z0PxoJ8V6MhVRf8ZWAoxivRLTJmN/vEh2zBt7pwAqA8uW+CIafb5GuG1xwW+OoSINLSa6TLkOOYf
zK0yUCfCV/Lg4T+RUOq/Ao1TBqnaESyBYPKHMewpjBJH6cDb5hy6KU8QsEU6oYKwykbk60tYEFwk
BPkvdFXD4psHHq+eDEdglPwVUhPHD9nGyBu6IJFVzeH78nYRpzMVDaqn/E8xkzkjz6mOvfy5Drhk
4RbuSXKfninmIVZbhzRnapYmXBOygLn9k9jOtf+bkQEc3xppXrvyqNhlisa85ww6+FPw4zI8d80L
qqTTkxGCcKWOqS8F2lHDg8fZZLf9lYygZrc5bw6LV8sUEhQon/RmIIlaWCpdVqmt9opDQKaW82Pm
JNcaQl3FpJBITiR7i7Stj1sQhGnAv10mdYX0gTpCJvqRoP1HhfnPGgiI3FJVm30/FtQyfyDD78tx
11l/KIfJgKGuznT0m2L1pbCPrBHF4KfxUoeqCbDajJOcXkn74C9q9mEplAPhYh2M+NsTTTgszHks
SDK+8zMqlb8IiboO2OBnI2QqHI5IbKcjOo5eUkY8lOi+oyoT4jwm8DA16UajEBMSR9MSixQ8CI+6
3NXfISfLwsiWul8Ed3mh7ydJ8+ZkK8jisB8BVXa8YXL6zezerKSv4pe74eqcfTgHbfIAZkxw1vvS
c/2xnr12kGsInxnk5gXNbaCdA4SO+AqkFp5iM2txYgRbFaixcQ2bAJaLC0gnD/YP5fWQKVagz45i
3KWyCffM8o2IlEUbfUxRKuqhjI9mgpA0kUGD5oXRiShevVrf2JYYo2Oa1xduv/VikeqTo8ILLCXd
0El8go+2j6SGyF9UG7VE1tcs9lP6hS4cFxhLNnzliB6Pwu23Yuyg/1H9FKLI5k0NC9BI5SneVNit
rNF+96GhVTj36uso3XzvPRdV3GQzWD8lNrK4vQlfRIwXU4L9W2mlDpU3vgewSQSHoJzsP2YYsen7
vPrUtLde8k4Vexr0wfSyOwKywMu+09LFc5ZCribM8nBwHMuTs+p4l1gFQsz6pB/fbN7K/2gL9pBy
dvqldJsy18KZymmmP7+ZPiibjizEij+qxGJ6FXdMFvwsGf3VDsn/2gfy4HyF7Z44sgFPy/K+6gL4
+N/Ihd5MUO2ySgLrbNS/gQAKgFN1NabiDDSbkfQ2GZo+fPPMQVyNJCEilGdlnFDFujNMcOaogD+p
0/dZIacoJbk0okJYz12tSm9PzuNwpAVH1OOcOuF07e9QnLU/9ny2KVy/lqxIbdruOJxfniK1JmTt
XNum75yrz3uREfnHJZVSz4EaAn1qgWSn9A6ZnDzX47Gzzzgb9eSL9F1fHyCt0V5nuiKMCfV148B0
OSqlcv9YK3sKbFoL4d6kM4mLLDOcvOlQkhRj5NrAcOau/Iw9PUdQecvJC/92ZgFh1iB4U756YN3G
ohkE0RcmKn9M0HtKJu+JmxDWhK6dNR48Nff9qFYLEsEhbLhwNiM8Y4bHycl3/umCVNsOfqiEHVaB
lk/VGmynuAAuQOwONNoSUcGSJiXlc7dXsqbjuw8L1e09qBdgyjQ/ao+shgvRtYJV97pi22Ym1yby
v4aYwjUEXGgzdIocMnlC4M/ifg/RyWuJz1CKrGLij1iDqvnPbMZGjTPTeE7hlfTBw8MgBVEdKqMs
XIu5RZindJjzyNiMt3GsierzSHrIB0BsnttEp2aED6eiyfsNvTf3+ktHRv1zY3y2LyNhoGyefBTA
1VVuAtKcAY8LcNfk00f2I2eQY7LM5IBtgxruMFi7I4A5DF7cUqgx3TyvTQp33LiHftWSTaoB0xfx
LETWz00mK88cA4XmYkXB+mQaS96jSW52zODf7dEBQeJR6c2InGXQAltJR142357dYBg3Zl//hfzq
pevF9jaoRWdYZlN4EN6goEG2pOiHiWGiBfwtqj3TPaHmUSE3MblqaAF/297Hokkbg3zP8dZCfZRJ
3vLoiv2BHook1VlQPhIQCU2IB6CnA4oUeEk+pRvvPWHzHkIPc/X41s/H4tp4ENeUeeBLr9bVzEya
2mxtI/sOu4191NCWNhP9O/mhK2k/SGxPTZdP1b+Bhc4izBGrsG8BRi7fQN0NBr/QcTAcba37jSuq
TNmgFSh5COO4fvu4IhxUmTxZwgaRhv33pR1lGX6rvdV8xH1SzxWqorLBCp3S1tcskRGQU7EPdMfT
gLjGKHFraM0KVfsf7xX3CW6RNabPWSHZDfZv7KKNN5SrHiGjGhcw89e9aSFilupybTITluhf8w0J
TSElE1mRuwyL4bTrrZhaJDjUpnIkF68v0avOxF7ClIRi9V54TEX7CHkD3d1RFJu11E68l8ULQEoW
vU4oYiPectiuiSE4gr/8bqjNgfYh7NH0mYlmcyELcCiZf88YGHoiuwPEjK12xmI8wlWUk03Z5/fT
4Dkd5NoH2ja+CShmGKSEz4jfi48QwhIsK+QxmCOCvtGqkSRVcEMdJGhMcJTSlt7lYtRPA1wwNysG
iC3cST+QUX9m0XlY6ufXnDRw+C5LkMk3sAYTujyyLwp7TcL9Ov4wWqlw4D8dFhHvMlh+kAINBfAA
pMkdRPMat3LysLKVVtgPKDB//xGJkAJikyncWBg1TN4ytXQ3MCudIWb2AxJfGzaAMkxpE1LAmscg
Tt0bJ/og6EIPXzmAC3mwbS0ozew2US7lG5hAvOj/DFNhjfGGDXZQwbMtgEyGWeyp0chc0mTROR7U
40M5q6xAW4WXjMV0C17oZ1+Ps2trrD7crnAUfE+liHzAQh3egkUu5/N4cpNcup01tZqq72nDERBk
VwfmFUoEDzrnfrj4tCjgASK85sG0adfdVWrbaGvQy58V+l632hTgFTIVOkFMrCsh1xxZGP9jNLFE
G/zF1Ck971n8Yt6f/8iRhuwIshgVsKeqG9o/KXp5m2mzm1xqQPyDdl1Otw+Q+ZAwpr5iDhutLJeZ
U5+CKqBbiRZYv8hzwGATO8f+CWG3PoEZrcMOHUzYoJAS4ZITCgnuBiEKgLJf3VfnMiS1LMa3qr9R
g2v7q288vslv0qDT0mdipDuJtSUNjnqLAgLei0u38EKMgnOg8/0dhXEt8nD1nZmXCz6Y8u6+luRr
KmiLL7z3LdTUI3nhGxdG3kXGCx8cCshXqaGadyh6/wl0VUWY8sUI46D1+fttaDLF7BMzSbVfqfBX
PHGb4QGtPnW6ZrnHFpt1cDpRvs31dcnFgFd5AEAKdp5ppNj8gQKF2Ek8yvsJPGPWxuL9rT1si59T
NUsEwbDznLVo6oITvvr427YuNMWk2cwJKfS8qHf6WEetUkWUInocrG8opNyeD9B4ZORvjY+bevMA
A0AoK5Ma5gPS4l9UAu5BWltIH4fIyPLhGfN3Q+3vHbDZ15cBuhnJtZnjhhKYP8LvhAMbnapORifc
aG9ihZwaEvoo21KCEBkNpmFNHvQ3uY4dt9v2ugKJxb1oZD+bG0Xklwh6nQwFemREPomox1I18pxy
jeRy/Y3aB31ff4Z9CZHfEHlJ4D1kM2I4A8wSB8evhJSE5jvtJttR7Qw6bL7Tvc48hzd/HpWCT2TD
vu3tcjVQNusUaeyXk70ZpDumbnt1HPqsRR0UPmcNUSjFJpXTa74pqBNS5qIpwr6868uWBvh+BiEW
sIq9zK75xrvaiiaDNzAGNV7LXT+pauljfygjTwgAoSrcOW/PgdVipSE7P8F/jYcob1AFsFOUkKM7
/jTZsqyLd97LOdkeq98wEzA1IOW3J+YOAKgoob2gMWL9hdKmGqIw69wMgQiu3Lru1GnopGvCbMcc
jHKgHovzcclGlKqrlC1pJUU1HqA+dKV4WIhgZlQ6a7QmrR+EeYg8NvU+pY4C6XxrMwDTqipS45vi
0hHXf/utrIJAdCls3+NsTsLvMR74oCcHYAsCJCR8SoNqDH6upu5B/BwGfWjvuYDqWFuuYGK3AWaS
WSGwKCEu+cen2IJ5Jqy3KJdBKKvzEFo4aOYykon4mYe3cTfK4qnLewB+t+iit77CTaoHRgjrijfU
fI+uZ6DFT39Y+Pm1jYos/xOYc2UzerMbvxmne+2LE1SMWiDRlLvxgYVe36jw2tZ3/SVZKP2Mio0t
WAB7KJf5wdjxCLSE3yJ9g47AJvtOGxhxk/qVf0kg9o5/6BKrnDnYqyz95mGxP7N+1EChsJi4/B3J
SGWnx0tE8qs/M8acAfR1JSnMI4HcOnne8VBKgrGEQbuNbgdxPt3GeM4xDn1KqN0QiMj3Fu4uNopR
BsxaLwMLxP+0tQn6ys8FB2hie5XM5GZ3ZvtZBI6G+CON3AR7UO9Quvjf63IVZIJvYbipaH/Qlyt2
vRCQIj3XlgYoVh+fjL3wtsD7tVzL5iC3u94edfNwrx/3U1UMe/xokEIT8Ept3/XYgG8h/wskbO1N
lo+uM/QxyY1ziY5pFZn7UfehH466iWuTIUMKpwluj34y4osAMnLKKusFOC4+U50AD6gStZ3TfXKO
gRvybnGG4pJZ4C7Dh+pwZf62zUKV7EFKI+4rAsvU8KqTjnAelfANQD29qSTBXkr2jRc4kOJwyWJp
MFv9Zkskf6HhcNUfgAUviGNvm8CCWijlAMOFqLFxJq+GDYc4RZ7LCNfvHj/Hv0519ldi2MuU7td8
/gIMvXIUAnRRCd+PtG9ZMNjcOiXZoSqxvFl3UI0GGdp1Y9l9o03QacoWPm8Hxgpi6ftRSsjcg3jT
YLnDy8RZACgp4TYDnF2TcndVc47XMzTdlcZH3gGG2R+Mtxxe+6Hs98tfYRcg6j+4xLWITm0SkbAB
ECTK5y8H0utlpuV87sI8cy2NTKxI2GHi+w/Hz/DyxL/qcuLGBQosJ5Oxb76vsraPVHNYvhsoanMX
tsVqQWQL7epbmkVB3fzPy8BRxZ/ZSF/vx2zCzp9s5UwBiRwznl9AfA7Mfd511yQ/+h3SCK9x45gM
xCfBTzgcFH1jPrSeFZ/uNTF+/ngD/sB4VpodLLlZ2txsMVAvVqHajjobkjStn0eFeLhms7yCE42s
njb6gmOs9VchbN3bxblujP182isq2l0cII+VBPJ2tL3GZzeQzTSgQO8dtZoc+MyTulBgUcZRfic+
7hZIAQPttzVbSsEu/wTONOf7LKirF29f4N8C191aWx/Vc9rESnxyrEUsLw0g+FC9Rhq3Jl/KeIGg
ZrPCvN9zRX3S1PVS9A5rTH4rz8O6FPSsFV9HqS6qNz9O0j7xt74fbJxJw6NSc4jLYzYjX0P7W6AV
ghC5oDWaPI16JTrBJGXZBjH/hthdmFCPbK7Y0iuT12idEp6VficrwF71pJ2O+kbmVKR/uxPokAFm
OubjukfqdUbZ9g/Qm1O8f3jJmz2EbkvtdOym34KkiFabspoIn5qT1JOaAi/xobbpuepylnANWQRE
I8Fa8JdX5WII5zcyMOtnYdbI+s28O5wobGdriW3IeY9iEjz1fE2rkGicqI2FkYEfTAX30OYW/4CN
Dx4SSAtNLACgprAvdF/lkX+kur2bG9Ii1n29Ks4mQQmLlkHfSkFZXnGHIssoc6rqdIN2o4XyIV9q
z3VFqGWUF1B8vfKq1ytu9Wxtk9kb1cN4pay9c+ChBCrSghP8U6gLUVa1Kx7qG3Tpx6rnCOnT7B42
nT2JwsVEPX8acFP1PfujSBiAMY7gCtj+LzCGt1VH8INR9gnb/i98NSW9cEn7soBhsN7Sf0VWJIAv
lT8dwNRdpY4MCe8HWqeYQrPC80ag3V1wIOcVoHjqR6g9AHdmJ/QN7mNKT+1f3NCcZPTpfoUvTZzS
DjkUUlEbO9DJZ0GeaP53m5cOMSbWgKTRYdRy1hMC20ov2IrigUDFLXkJR8dr2QPgdHz97oz36/Ov
4eHPx7oJIKpFostFqJnROoak01DuXw8d18IUZEwNKCrH4l9q8GfQbxsbAQIabrgjIk8YD9Au9Go7
wT9RQlPAvjlqkk5OKVYXIh+p1zPXgvX/hxN7nQg+Q4Xk5QHHRR0JuICbche494ewLRmaysaI9P2L
G2hxVALl//Yrz+vKndG4Bt9+zdWmrQnzieCdTfd4xZ24NaPtOuVN0ydlAUAfYFMmngXITNCB80l1
a11J8XB511MecAN+6s/4nYQGtyWBeBcBFIKIRxa6UpLJ/h2I32X4F0dH114+u6/VyIXbhYUjP3Em
DJAjNSekTnDVHx/DlXn/btyIlepW2kviR8FndJjFAffVMfMfuhN4BJLyhp01SsJrO3f0zhL8FQtW
1Qt/TmYQD97/u11O3eIFBoqkxRevTjyU/FDe4rX2zYlb2ia3EiseXuWncA39hz8J9Sat78uD8Krz
QKNCmGFVzqCfABJ6TndFJRhGn9FDGknV8AHfeSI/0ustcD2t9Z6MWAasHNSuHgqluqEre5YQ+ew8
rm30SlLt8d4BQahsL48cMJsGGnowwQKgURxr1wg9LNjvuYZ9yeQXHIbMntSVweWgftb7h9wca8jQ
W5fHaS7l09X5veZZonIZjT/c7Hku2jiH8Y+c+Plxn9sgJom5w8JT8zIoatlYj9sXHzt1wFITdfOy
A7l42oZ/d6Tnc7UndWNRdxSpjdGZc/Mwb/t2DWGti+XEB/geZLR8chYXBq9lskznabRDQi8GGaj0
1Hvn0GiZXtqZ3HT0ylO0tB2G3LPtjEht4J4ZW9xSEv8O9MTGoedrv2YSxnyPElpWdF901vrbKpXN
KuBBjTl1XZ8k+AuGxWvFX9Nyfj4f3yseLK8RfFgr48PZXPOeVcXNntxtuU/93rYT9Mt4PEIv+wyf
6lYpHVeahj/QxtWqt33mdEYz8G/5i7lEym5HpwxAGRYt2W5cBmtPOF1gFFwIQdaqJ2AbgAAOdImc
YYNGCm3RdM+QoHxRyHv3UlUTGIDna5AxwxqrlbO1q7m+MqJG/AdxjTOUH7M218LoCDBgnWvShYNP
i47ZFhc0NCPUVN6I1jmKpLHFZW+YGIUqDC8rallv7OByF/X7dcPy5F2TBQT3aZVcaIyaFescTvp3
fnVF4ga4qXqtP8b0JvXMPyA11tnVhES73935LZj3YxP2jdnROtrfPQh/39pLqrocc0hslulV9h17
3PfHGt+xnUn3Vo0WVybM2d3gmnFuTmUNTn1OlfL1W6p6LkY354GDB8Fk2Rry6+uOa2xQuWUAMkRe
KA35iFQXqiQSCi9cZ+/pT5CI8HDO+Qzth68AqH3eKKz8bfsH94Do4YxGR7KYztHvFIn8/2wCeYbk
bFRcne5XZAUvJuP4P1JwjBMa1JE0I9tYPgWj4+aughPeqQefKvSM61H3ygLOgfvvVdKg3ik3EShl
4+kE8XPO3KmxenflhS0Zc4nzHP+bCgCRNiDzFHzsOKShKxR7UHbW+DWjQ8FTAY6F0xMsR6cXERkV
lcBBUtiWpy+gGGWjq7GNSZOqnEuxl5/FLDmpYeTdCqJTW9fHsqKnlla3hcbsVlcAOATpMdi9US8A
evOFj4v42p2+ce3MorMwyYaPp8u9zFCfDpFRZvz0kBgzycGeG1VUYNzQiM+5UXr0YZ/QHtKUO53Q
WGsoF5Ew+DotPOms7Rliq1G3wUF6cPZeFfcAo5jx74qrcld2PH4zwEkO/Xo/AmjYp5ARNWPqETR2
R9lIjndn5Zc7KeRw01tdIN8RjxfDoUK4fK6hCdbRpZh/9TPltP6uhEwnAvFyhLmHVzyZfOP465nx
k3QCkyVANhNaiP/nlFxAeZmYmLmd/NBJ93Se6kG9faQN+rF7jtQXiNs+oGvhq8NAdjn8I2LZDqqE
7obfP8UlRGwjZ7L/X4IU5HdPUMndiOfkZAutzHtG1PwROo+KIL/vKoDXozMhWTsUh0gPLduVw2fQ
ln9LbEZIXJsj5oN+wEacODYHWzT39ZkHRnvlHAy+L/6PzQOMqVC/TQwxM9A2h2F4QxMmUBD9yT3I
70lI/m34EDDSz10uXDBmB39r3gIeBS7SFGun8FSohvJAmWNlCp/1t9xRNVrlXvj1tEUc4Jpbcnbd
tkFLNj71EQlenv8+dv24eKEew9FvKcoo3nBXzY39QF51cPqQUngeHmJaxBnwa42UR3Q9Fi1P/Lsz
dhVEoc3acdwW8nN/E8uOEZV6e2AiZXKWfKL3Xf3c12PiZmVfDKXUwUOQUYsgdlK3PxZwH5DyuCaP
QxStsYQRACty8M54FIS8Ycl2q48iIQUtKszAPIjcnaXfIg/U5Kp+asdmXbznBaFVdFywf7uT8mvd
jpQhXzQUkVKYMgG4iBGmhwj4GFVM56GZvczsNLedEQcihbf5DxgdL+JctlRu6UGUKF776AcAU38T
g69xoS0OWSm3e+TDvDQ+iGUf/Mxr7dbx/UlG7TvCIRqtW4YLKzgvktMRUQJ+1hu8ZJ6yRRiihyf4
ewjeTie+F1smcgVr8wir7naq6fLUxoYT71HHTWWabL5uexCqdsOODvBKJSX33HmMuCRq7YW9r/yq
AWvgcAfQ3n8jMVUvX3gx49XXCyu0ojWoAydATiqukjwCs54tr7zqeXOMEqyArkikzr/wqIya9LLr
4MzegPd/NnmaVVaS7KHAUApioOQ+1Q6wxF7jThG4cHjUvJAJa8EIbX8B5MFblURnQIBmSuQFbYMN
ArS0X2LhMXKNhCCCI+CuEDcAcJ61zQSB/6d0hplAWFXAbi4XbzzaQtla+taWdwsUQWRRw7ZdZjAI
KYGuqiUcOITy/zgvZCaFhBuSxO8iGfJ5ntZG+EothIf3t9dwYu9HN4V8ZwVx+GcQ3gY4vWLIQ/NC
oDuMk4N3Oc6lKaob4Vx8/hdu68CIrWeDrmMwW5ncOwwSQRlrpUR6jIrQMyh4UvmxbwmjGaz66urb
ZmF+gLgCEiB8FigLLsriZp3lbPlkXSn5bjjhR7XvIu5lotadCDoDBBVum3kQgiEHZ+RdeaFh135p
CEAh5EOCUvXxXkF0jmIqFSkDtJURiyaXWJN1C3wCvX81mawMLGxLpy4a2jZJldFp2fOs0gzghB4O
1KN73PMRv9lwdamYZz5axNuVijdqlWKjuieseRl+WhiQVzpNPu6LKlaxA0t4e2C0l5T873YvkPiG
ow0DkmZT4yY2zS4xi+2kTL8tGwVIH1dxsu5igX8MWsmakfrbsBT+8oBnR/nzWmUIdG8Q4nzZp0dD
QmR01yglFvy14AedUZXXwYbsJ3qgSvF8AABEyIYI3dF2pj3BZDfb8HIQ7Yltjw7k8UNRlqIh6pgH
fzLfc8Nmrgdgb6DbwvTC+VttCoN20ncmnowTTOv/C7X4AelGnqCdYeqsh6ZvARpra8pzuGxzFZW0
lkLqycQRNhgfIeLnfv060AeLrqK8hCCSIP7RSPTJBJz/XD+LM+6R/ylO/1NraNUI7/MQ3qKm4sca
RD9S9ftbxV8YTfOk+rudEiOMt4+FWUQLc6jLMrWLTj1XyPRhZt7dDoGUebM8aWbg1LZIG9wcnxn/
J6cnD7NMGRZ9gSNrMRDVomMMCXNA8PsgOmkex8oS+QXqK90ctgWWgTB/XcaS+H2u02joiWnD88Gk
RiGocJxaSMcRuYLeFH4GNhkHV+xPaDbALCgRs/WOXZaBk69JKLBfk5J3oQMSJKR0TUVXGNa3C8pL
cgF/p5CLY9qc70n5k3qWqac4+rfV0ZhY+T2h3q8l8Pu92CfLbjZ526dJBLZsGZi89amaBRxM3Rr4
ca3otRRUIrsgSOZXJZ3tSxVHwxF5jQQB302AaSjSzIjtF0ra+6EnZnBe5uJqECuSiLpZJgtaJxo2
AnrBpYjZsLGD/PqsRdofBIYPAjZ24eibOlLaCJE87zz+Iz7lE5ZwGErZOqP4tBLkwJOaZ6G3jAGB
NszF2zZQl5xA4mx08rOWWRWuIv3fZteOk78efEfTPOGALkurRt2Ik+K7GfxMi0Dw8QvpUcJWxQml
+ndhBxmqGm1YpryZAC1Ycz+I59UxpXRzs3Kxf2Q6c0iFPAxJsKOyMH5q8D+kcC885TSE9/gVTfds
I/oZm5RZa2otKY3S84LJtl2p5hZmWQSzJ6E4Sjk0DN31/BJHQFlsCxEdSnOxELF55pIVJjQdnuuC
7zzF3ypV+AjCpQ9obFJOPPWJRGW44LUZw/vYB6sj0Q5+jXf+jIk8OqcB6hC/gu+hrArzVPkpbSQt
BFa1EnL7mtkkTdkL8BURycdkoA9YuQyqbwAg93GZdOMZSrmPq8lg/pbdIe2+J5eg1zkAnTRj+7Ee
Bz6JbhTFz5uV8P3YSz0CpGN5KhuaO62/wMRW7rrqG/Q8F0GbauezWo0xf1T85x2leISX672VFMnO
qMR+p78kYBk8Qk23uY42yUFCxDhhMjRIy0Zv+elgoz0C0vRxlNksnUo/Om3XRXG5UL7NjMAlxMlR
bCMcCo5mVW9rEi4At6eSyarkOlwoyJaIS50vVed8YQJhrLCFkk2hwfZKgGd0k8XRnSV16RHTZmPG
2a9/z/kzELvPzubiFYXv5dhHvpIV6hqwnjNkU8j5BuFH41Xz/fgi4k4XyM6MIJpAV/xwaGcSUa1P
tFCr8v2MqMbT/Y6nFKhxJaQzk/G+SWz0IGGJE8jJl6fI7h+DXBrd5ZNmmQFkjA0EKftK/qXWC1PZ
ZTbOwGdf1IbBaLXraJiG/Lu9GrL+VjOJeycP+GUjkx/0lUjt4eBjz/UCBG6QjUmSm8Tpo18aEFGC
vM+Fwb/bzCUzIs9WhijmBpQwai29I9ylvBqdwLj/5Nrvl5HmcgFHS8+L4C1QqViEgTCuZehOhEh0
KoUTxWe9oj89yj0SNAl6ddXdTo7ShmM9U+yw+edo/DlsEO8IbqU31AZ67rrmZLqkWlFyfzO8Pq/w
iDKKJUsVyZ+6xNr253cwv7cJkwqc0WdZX3Jh9Ph3ecGpRUQ5xsARV0U3v6Za+j9oINZq/271keDx
8Yp0WAKXI6DhQB50iQCAwkLYhCxqRMLyxd9xL5X17Z5sAQA76TeD1UL/jjT7hr2UbeTcoCThMSU6
a9RAR4sDbzsIoNDXxxYUFSZvH8zd2k+j0LSWSwh4cz9q6uMaQ0p/23h58Ttpw2iIoEaXnzTHLdq0
OEBZxwgZpcPvO74Wdaj6IlUHY37UHJaarsATCOtzqhZPHm+t0i9jFWkBTNXXJNLQ+8ZNEc4eyurm
+wtMpJVMaMQdDbvrQko+NceIvlOEkUuGW29CrD6MwSW8dLBU6Y/5NDYHSXdIol1AFrDfxlTZutI9
mT009Xp7XTiXFSgk8+AL2tPiks2RP1njajiK50IySclIvNDMsmj1yDdH5xN9rIfO6s6GBzvg7WzK
L9Y6GK0sN2vnhyI7aIyVHftMflR7duMnMr5Ym84whjr5CAgc5KabgVE/Il/oamdeffxEXJIeCqNr
+R8NVSxYn1L8GkfGAOrrr8whMa+cuUENM1G59Xp0/X9SrWKiSlG/lqQvLw5k2X1eqYdWIgpKk2og
Hij1a3n1Pm/xhqBusfT+7ORkLbzCnNxSz4o/W4tgPTqE2xQ5Hs5ARb7VrAgnuiUdHgQiecD0Bal+
QPrlBJPqLyWFor05quicvkLQfsahp4pc/yHVoPsTpRkIxbjRjJYSamNvxA6rrsOzE+7D4XRkzGBS
ZnwZKBsw4XGpX4n73fJOq9z+JqMzPZvqvVzQ2+Vmmd1jUhjvudlYeaV7mDx4qSBa/PKPxlLJRTo6
CWy0cW1OTA0k7U4PyzLUvhYVwssUKl9Q4qeSjHrKyEvJ/TRbLhlxOZnGm4d9azMn++fRzdz+81H6
ivyvVEusuv/2HplErWXSyQfHdgKSjoAMQfuREXj4NCbkvao23M1mpqH9fBoTeVVyfUNzm5UGHCDh
0Q4Q7KxaEoplKoNHqv4twCQZQOp+LXLUlAcECsklV7RT6ttMjvWA5m/QeO0eCvtjSZuIGptQO4x8
Vs58uoaKRGQ+4jgedJ2x1PHahBTTqLaIWz/2vHrZwQieFgHRfUhOorNi5HLaJTAm87puSMBBgdoG
oH9Q5y8mpti0nFWQzuyef93aWM58qbJfRrFCkvi4SZ+UneC7nf1zko8AFMqQebwRWtFJba3qKiN6
wC73E1T7QJaHsGFx5vWF6cd6x0ZzlV3mP694/zebjcUdO6gjpcMuzkaZBvePCB9wWLVZezlJd8VZ
3mp38ieS39zqw/VEseIUJtgbwPVuoFbwMxg59t2DToEMrjSiHwvsRq9siMMxV7viIzWFG38fDxx8
PwkY4BFnbmp10JlctA+8YXb+PBB3bs+Iu7KMxyayiMQOqDSmzRkhOkTxvMshrqrdyNcr6mAKF1Oj
cD4vBmPMzoa98cT7PI+JIeb9/peDvLChaqjHyxozkZvRqL9I5zv0aQxmfwHtmafqWiCIPhk8Lu4D
1sBkHqMjXbKdaSLpsDplmmKfs/6ENPPa9tCfcRe1yEP6aWVY4+kN4cJxjB56WMMrkJb23BmBUVZY
WL4Xnllf0FYxL5TTFI5gAD/XtkCBTasKafewmvrispmHEgCfVEF6XsHvA812RW7/M9O6koilG0ZW
I5P0iHQUnxbQPBMm3YuRIhSctLyE654Gs3sW81q3hPZC1C8nVCodn4voXTKLPCckcaHoGU/ORJtf
iOsz7C3zSZVV0ZzG3CYmL6+MF1A7AaAczNd+W9TPWJTPbu9gmxOC/Rqlry/8Ls32mb04tIT8/6WP
Zp/oyJtPztHzcUugwoyjtNTIE/vJNQ0oc3WVwmQJq2e7I2NgFt83CKx4KC9y+qwUVXEmMEfaEWeb
SzmQNwlEOiIKoIHk1deVL+UQiMOOD/c6CBe26HpHx0LmVyLy7XovlAz4KIrpVXynG/dDGMrkNV0z
rGSedkirA1hfEc3FG1WTkItbXtXUNh+6NiJPwqQcd6k+n6b0mNxQSP/gKVqFg6BskVokkZck7rKu
L67KNFrDP8Q7av5P6o61z7y2keH8jGaM4NwivD0n3yU9ojRhIboVD6c38KMuq1l/o1Zkm5I5ToOI
li7gQgY7v4m1Bt1a52/vgjYyb+G2CffoSppxxrg73qF87SBa0C1VS9AmGIjHqSsoyGpdCwPJAgxm
EzS2+0AKnv+PQuvssHVrvfIxI76LG1F9QmglCxPmo3PHE80oBCLot2b3n5nI0qjOYKLRpVt2K93p
yGBSq4EOKH32kaTw8a7lEc3kDsyb3KNECtcR0B9rLFphC7LNfLD3DUYxX1fUCK2TsmVSTu3C+eUS
ZB3Ib3YUqjLSSg1LMoMsuWE4q1N6JE9WcjvU93PJf/G5or4iNdv2uQBlctNdEKh4ERCbIZOCuxhB
V5d33oYrb0OrGYdm8pdbREgoN7zfMK/nvvqAcQVEQVMsO7haYdcZ/S0IOIbEqSaRjYeOlak7wzy/
Zt+zTygEZ69eVTW7Zta6PGG+Z0cjHR5v9Wo+8jYomPGMHux2UwIEAs00RrT1WQlLN2XT2lZ2Wm2H
KYWuzskx7ig/PHsQbs6I2wJ9dTTHtYAKFWnQJhBAIkSH2VqsZV+clV8FKUorJbnlmnr0KJqjGs5K
5bojNNpjHUVsJN2DHVdMgeDbKrQKsGuM43W2Bwze8qZHQofnwETM8LK9o9T4ZTcE1zSZ+sF/LvKb
rpTFMIzA1VMAq5kzP7w8Lyq+FZIOZBGby6PSSHi3TwhQlHQJvowOLY1tt6mLXcUQOK/YnJ3x3Aet
J4KlC9oCTbGs5hz5jDtxWg05vumkTELEznpuqdSbOOadmyxSzA5eCbWjC2AV6+r2goHwyzHMNLpO
H9lbMpnqmdWmwAlzlkNGD2ztYC63c5U70H1WwJPXPNd6kitE0BPdTYftndK8lUuK0jqfE82J/TTo
YjjX0F4ubZ6NJHMCo0bLn8lvK+mMw1q4TwXK3t1nMB7nF3T17di2WXQPUya3Ljgui1EVJ90/3Zly
eASiUTG1h0GqCXXjvAj5liSApMqtLiXQVsNxV6tssubqQSVLVObtm5u9h6FCuae0w7r7Da1TCmzr
oVF7wnbAdYytSXVypx4xRqyjWGimyqNPo0p48o5LMaCDKjRCt0irvRNcDxkXq7YzrC4kTLTgKWuK
e6oPxli/ihj/bGNUFvVa5H9uwqwDMnT5kC6YfT0PoBIKytiprs29776ZtHj5mBwJ+yo0dV5NHV/2
6NpWMhhBE2SGr7pa96COg8oYeeqVuzXLjJ848WGMPMe36LsMc1RFbZRIJS5l2gUr14TbCeeldwtO
xBr0JhxuZBUH005bmR7DjvPKwE3M47gGu22ydMfJYs8XspLJ+fgLHB2IhAl2D0uDVlx4azEwjn0Z
sx7YKakjzsY3z0SF89rpXX0w8KxdJhbnwrZn10AaQ1v8TmUTZ+dWCXCGFXg3P5v1yekRa8goUBva
ypxJWiPc9EGq8Pxm/p8QMAKHnZkLCgCQv4zpO3yFa3f4iIRhg7CCy3bWzRNNBEFkPVLqJfuY3NTJ
qSUPEEZ/WM9J8JrZsx/dUPgHziMkLGj5wiBcqTGROXb8vjg1ndqd7lKZbPAsPjd/FCtPxz0d9jI8
NhUPHMUV+i2blMaFhJg1flq7wVHlVATWjOVj0oN5xLJCPRjcBzkPYepEee1NmYF+vCwOaNwuB38r
y4TO0jrdhOwo3FjHqmxm9qzo8Krpp+qsPQfeiTEeYloteyXS66vY6I2gSxzrSGDsMOrEqKrc7kHt
mETYt2VMGT6yX9jAqT0dgICrzV0pC3gJ+YoABfyXe70C+9bGNnqY2qoylVqdxMSZtG27ZdTEvFaF
E1Yd0/yyYZJGrC489FwJz2jZpIXfoDbUOFgzluVRUz1QQOtn+N/n0NmI1gRnWDBryw0jAPZq/U5u
tTnIkWhBuvcBBgAOsOCwIgIf9x3t/0gYB09d/ey0FrCyEpfATr5jO/TEDlH2gkrIHkPhNCYtDdst
XaLP9rt46THOF3o/S4tLiNdtLr4qL3911Jj8+yCbp34wtV7QQ+RI0dtdgwe3aNyZyOPmH12zOREt
xudWZJnPFQxGfA2NoQR+oLVO3X3T2eggbaamqswgDtJcpQdhAwn5b0CtBd1ihexziJXVuXQUP4k9
83UZZHOiABf4GckLaYFsmlgTxGfOZgw0NYXRlcGOFZzlYDXym/davNJ1Y39Jv04flP9kIB2j6lB5
50kdzlvZN42WDMXnQu+TexGzNflIdC2gzxAj3g7YFUEltKk+SVQJr8RT313B5D9D/HM3Hho+85fH
erCEmhcL1ThqB2dShZ57jqrXAfWlNEdk92294AJ2ZeVfaXp60Rdrui03ql6nvSOGkGVYJlJANA56
ps9vRtOIOQ4cfWM1RHzp6DxqFyT29IunMu+KjLJ+z2Ws/x8JWWWGpCVCgigXUc8s6mE0r5thjr88
1qWdRdzkmCQWTQaNWQo1qqY2ETVVTEFO08Bb6b0VN9fYfZtGbqA4Q/JrWZgk6ZgjAyWAuvfiRdF2
lw7IdCVeWIl6JgawuU3/6sbQRbQTTe1TZhDvCj3CBqUMnnqzERvgeHIuArtrhtq/psKu4CqA0Tbn
OwozbBo9YGydmQza5Q/Ex8YQxGp2R6JxtqtiN1JDNA2m6P5kC/ggrIaLmXyMH8elT6/swArZffqr
ZnrXpjMY/Yg6Gh87+R8KyGKxwugDHoi29o682YhfhMNhyYGrpIrKCTHYVMR/ijcu1vZfoCQWmuff
clNr8JKOGrQGOJK7dUgDL0uBaUCUn0j12iQ2piFfuPkxifpnXcgKbb3cd+UF9ApS9ykAdkzTSSLA
BsUJUc+iOikr1rLFykzsuxA0zJtdseunMqZsQ/7BRJ8A5P/r+CvobN3JASWNU3y/cNozxL620zUV
bPQyq+au5F9iMT/ubVNWZADSuN/ZDHOjtdeQ9l/byqg166TeQ92nC2+pvkgTh5QURHXjVsy+ABA9
MB8nVFO9X3N2OpafWJpbswWsKOu9w6lFhDHFwRRicaXnvilJ//eJ+Eo7w4+ezushwTIz/UIdmE3w
cz8jdd4RHniAZKVYZKXV700/diCr3oQgKP1Wxo3uixZ7STJl/obAeycwFDv8JnoHx8EMroxHUTTN
x2+6P+/LVZxkNMD0lo8UJg+u/0ry6aisD83Ea5tcK6zc4ZLbv55MUAF9spcAcgTcqqGOstkvmLR2
1s0lf6mMb9VYOc/xjFPDiBA50DHfoLipPh6Mx1zQrkq+bccAp4Ti+0FwIJY863JRzqKzRC/eqxJf
eVIvhs4QjzPhkmTmz4v7cDQlgZ2pKjz+rgnnO4LLiX5mXYGdJhb6SD6K0f8aElCywcYYze942mou
ktdq2GHWxnxBI4nF5wITDbBcTj4ACBClPuUIdo5wSmrVsccRFmCs9H8vg7b3Vxb8px8YMDi3TLeQ
TQIlrMS3E7t7DBTM4MdLdL2aQGFCFHdMCAuBin8iVBKacMx6BaXNtGH51QeeQZVAOkGEHiXi/8Nm
NoJVI4NiYh5fFken/seAzsEtizL3nBXhpowB34MazB4UnHl0hmNt3OnbM8k4S2JrddFTUZa0uW42
n8WrEi2PSVeoiK2zBWLmFTSU+3L9OwSEq9y8H1ihxdOfJElGGBkqcQUPxqpvWNFl5+f3jaZimIhq
pw8WU7TTO4PfXdIdM88oTMtnND7rxGex9Sc7guOJGoK11sWWCDucgnY8GC+km98ZKCrZhu9kheVs
HfiymR1i2cquqTinsn/Mw+07TrmtfgLstOQMwZxBdszEHbvVnMmHgF/UIOpL6JRhaxPIB6BGdPev
zAiiInh9swsjOzc+cKPc7tTQDjK41KP5g6D2VOR8TZrljLjNSfzHxQeAF/pHzjzerwycBb7uB/bz
R5pH16hwfsnnaujnK7RS5kalnkonu2MpoAVJRdftCrPxFth0PJiXWNqrL+44KzZu5Fk91p0gU4bL
Sc0FJ2Bz2uaEbZlGUS5hrnSF9V+L1hx1EG/wOUVgxrzVS4azvu+syopZIAtBrF8LOsBIvgsM0pdE
SdJSSJwt6zNCrFhBu6iHolXHhSqCPTe9MZYVqN3OArvX5/Cq8U3ELUlOVP67BHDvBwuTEc/83uX4
M/OA6k4urucJ92MKBvOR97T6c3ty3c82EkZv6k/vCvK5lkl6KtG4Y+9DSVjJAilulHqJ9UaujtVO
iZKfQ5UozRbiOPeaMd+FA7CTNeoXtZkmC9eaulaUfYqRvX+Udb4vAg79wBo1T0SQ96PFq9+aIeP7
Z8YZVr09SMzAaAq55Y61BwiLgvfBUIjQkClrPieFfhk=
`pragma protect end_protected
