// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
WOYYpXv5VLKXxZJ/ix6VX7UUuzlwmCGdeECc5e+PO/a0rq/n7V4+/X/4nwhsDcJ0bibSa5tQVVDp
tkUYXHXzj0zKabNY0QvTlXtvRCXDEz96/I5gSkAYnht0Gp0uD9GaQyea2W1LILzrBYmwqycDZg04
O1cwM1lHiYeuhlhkhzgeGx9rB6NCC1wM1/4fkt44rOqBHnO/bMWEJtqcxc7N+lc57IgeduGaZjak
oxAdVUL/hXRFwiv2Z3Ln5hcaTdNpHQcsKgq5fZ1mshePxS5zcYRGMdni3FT9zJr3dFkoe5LF6VFq
uE0tI0rngouFKZ5Sf/jAifn11/73sAQwWx0uNA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 58256)
Vih+HeDQXN8Rf4hoyuA2v6YVc5VxREKcP0kVRwOUFc5k/RGfJ1WgOmDUCepCJSacZqrRo66ckj7I
vHwF2hLd3Ybe2geDHCEtjOQAzP+4JF6DNdeEYqfzU4+HeEtAF0MEY23DB2iKT8AlPnu4qfkw9NhC
Cb+lJb7qEg4UReG26KpOT2K+n+rVX0Pk3le9PjQKJ79nzOKoLtrUfZ1hOB85Sl3MXnawsFO9xtbf
RtxYGcg/wY0xrOkp8wmZPS9LY+62OOHnW/aj5WP0D51c5kYMq/hhqcQL4JXdGKRp+YV27CW+gaWR
ipziln+6RgYNc2uQyjmdHDb1tAcTA89qrIwJqIUVKNN6cHs7McD1UPG1PgkF/uscvKv3Q+OQxBKO
0LSZtbqMaf2yeKhpjidMXc0h0YsKHB90JPuWSeCixxVoIFlkIn59VOh732AxX/5FMW9a/XK6necl
caAOslm25cOZTVzDwSHU+pzhuv5CrG4K/Cab8COkM5EanTz4jvyFCuCfJzdtFogJsQ18mLNIiix0
TQ1bD6UcDFrxYeedEm4IdwlZqYt/t5VX8OH2ZXFv/6Kgm174cVnUI0eRYlXN1p8xucKmbfIFsPCo
E9rOo4k7LRnfq4CXmDhdsur+/6UswCCVlbtVKAbPIkPKl4iVD/g2llM3PnECF7oYRv9K6mU9rEV1
keYyXZh0ADntgxLcgeoc3iES6SwSg7BNi1KuOvADInlslIoKKP91VmA4tUtEo1bdzL7wFIo3tXEt
PFkJ/E3eRJKdP+W0BT6omncesHkUlGKPPKHD20puaQqkmxIGsABm1h513tDpC/848+3PUc+oKEAX
bImMoRrIPkVHJrh6WBsRqoyRQFeOalIUDfwe62bpfs0W1a9pH+X+jio487f7JvTbrXbnhravrMnh
fte2qusLFrAH4x0MCTQPVVyMTkYwR44rOK6s6INmbJqzB61xKQDxdxkEC2YFLywSV3RazteWd1bA
4A/pgMUD+aGMm6vu0tYfMaxSqCyjn45BynGauOCWTeM6QVoPEhjaT+cFTzSA9haGnMi+ruNixJ5D
kYnBY1o387aqNWebzZDPxjZD3gwQruErvaN6mKehgb7yUoQ3IHRuZXzjMFNxai7oQHh2TwKhrZFM
nQI+aHSPypkxzDekcMaWuh0QpTia+1nZKfLYq8a5qJKxuvR2uDuv4j8XDdE8HTQQlvlAggwVINhi
J/mnlpBucQiGg4xny21XPYiWPH9zEumhbORLu0SudX1mebMIfVj7ax8JA/uzgBrJLpsRwB3KsU+K
NW2npS5uj2McTruVkWnigg3X/n13FadncGMLDlLHEMPzcDl2dxzoEHpX2LDsrFw2C0Yx8DkvTY6q
8kzFfpZKw5Yg39rGrXP1kABwjm5ohiwHVf/X5BTNvSsgspDGkqWjlUNqLdccXfLqt4e5rH/PfEJ/
VBR+RQd22gVHaI9/8RIX6sLCRpBTNCwx0U/fPK+MUKGYPuEovwDaQxxYp55IrhhvnC+LSYiY6v2p
6t/cvbeQAbydPb22YQzCN8oYffuv2qcnD3Bf0qwhbqYpX644UdZ5M4ophu7P0UtiprK87dMqeMuM
bHCvBl3FKNFhdz4C/dkNvpcWeAcqdtwIaGM3UcEFBsTDjDlwAMf6KMlm2zZxTQmZNGUKd4JNITiF
Mj3SjzTpvXvOpis+DaniQFqdTIxMD/gZzSjZaZR+uTrp6M6AVW//wXC37zmqqXzFehLv4cMCTC9s
zK6xYWS86juu3lr8I3a51Pp1VYIK1BRaXWR4qsY4Ni9be32xBq4nb/t6b8RdvEN90dxfUZNy8/BZ
drkGVw/9cFtc9OUZe+V1vETa0HJ6mPafBNBG+c0+TUxGn4KwgLg/qBljfNCRdUKbBNcToWsaRW43
5E1cSG2YPDTxI/MO5OHm8PgS/846ytv4mifpBa2FKVEqSt97Bd/6o5uEV5yp91Fh3NVM9D2FqSBC
XzqxP4IGfKzYGiBecS2s4MDsHUxQIKupnJwkNXSy7tANzc/qGWF+yLoYzylRHwdZwJOrLtp2bS/n
igFzJHXMF6Ot3i1fZ3mnLkYxXkGMby4/srL0nnd2h9rg0BGfIWWiolFLCMGYK2VLKGh/K47JDDBr
URngsVPlFB8g0UGs1tHoE4xovbKMQUyR2MjbFFxiRXd6KQpD9h/CiLLoCN0tbi5lcnJ6s55C1fia
TMpcFxEs3jibLoGILSi5ZebYiBYjDhcRDw371bjIYKdAmIy91ACcBh+w9wV0WdKsBWA9sEIC554v
PBEfZnI+2aCpwJaL70a16eSFkO8Hj2l8xSG0wUOI7ckW0LG4vi6XG76Nh7jHyJzeCI2IvRZxEgYA
wEL2cx+hq5EIrT1tBejXQNffHhWRf3QLz+FGZu0C8ofIVLkm0v+IMikKvs9TRULKCKSI6D3mPnsk
pAF5Mu8XAkhBD2jFpZBeTb936qKvKwUTtsGZt/tnRFml2kZYGUNxO9dOLgvp66qlyEobWN7lxnTw
gHTx9AzUTf9QxfdIvVw4yEwijseEZgmQCJgHKQElh4ojrP8zLGGl7uSYcIrXoqS2j0NYo0zVO6ns
uERri6W7Sb+dVjgDx4XhpJEL8izXEx/IcT3TcmflXVjGXTDPn7kYfuzDNDfCN3dyt0o4bIuWjYHk
9HWDbv/ixv/TmtZ/jeI+DS87mkU+kKz3vUtWPUR6wCtrhCEjyvSfEalNjpsIe3OB4advSC0iVWAK
wp9NNOMe30oCKt4zyPAOV6tyK4EcHh5wj1cHDjGC/YMMknYqWCNxiYZMCIy1AwxcMegBmKynYuQn
5+SEJDvx3uj7DsCIFDfFnMxHtatdfjWmqlu8xBnLYTNW5Y74i0P8EQzd0pnlMZxwhkUcPK3V3WLv
FeFjQr8PACTIHKltZh9CbDht9NL4lGthB+G19gflnElLkDezg+GIw88VZCxuKRZjRcAqgkHLNI+/
78z0+Pv/eHZuKB4uOokgS5ohx3ZIVEhQkQBevPcMNMI2Tu6R+eKEunoYPgzoJGO2t0mAiEq5WEX1
JYyS0cmI/KZQXLNZmOr3ORLxaK0UpvJ0lSX2DH9ROgpTNY5wgJd3Jbt9OluZ4E7/rBrR5/P7AzUG
oa/XI3/clKKrUUNHB50mThxU9BZ7RZaqVfXBq9l4ChWc6+L32aRH7QRzfFHDZeG2QSWH8KOV+Dtt
evxueAkuxc+gAvev2T14E1XBh7os88Vf+eKTnHcEOV7ZtUV4BlpCdPxFPepxRAtq3G+1dhbZgytG
XKMkhlkSqYFf11pYNPl/w3iEN5LrvG3PcC8c8+2A1ENTsShZmJn9J5eQq9qeu75/mgJxsvIOXFsM
Cv/YyIJfIRVKVmnozPJ9aXZxsgTbKMj5fBxS0rCrFgoFe90df8lO0vezVcuXuMx+0Ho483oc1pBn
qXyEEJNlMV4NW+nqp1vufxcDZP3204E/Q9Oqtlqk2qXsC6mmxZOsunJt1OeQ8d6XO0JgteZq1UwN
+3DJjp3AqsGpOurpFhQvP7bFh9sOmd4uly/V+8IWaMyLPTXgpqiuozFSsGmE5Cb5XYYRAjXkjrF8
yv9zhrTVoPhuXFzrM9ZRFPefkndZ42+sIay/Buu0FalS4mWhaJK8ougN+monZR0mrFFFdguB+t2z
S6yJe8hniG80+gzyP1kJOeOqjc+dFIMGNQuhEBb+BY/Ayyhn2Osil2ftlil5VYS/nO7X3bWyX+3g
JjkkxVP+dxzUg51pvMmSin8aAghSyJcZEkx7Dztp7yQtNYFvf1cUjVACWjrc0aM6II41+hT6mD9J
jGo36eV/R8oboLHnVFOmwLFbNDuXTyQe5tgmmv0Fe+hJ97qpjHczoVLIRjOYQBJCKc4f/ggVr02z
uxoXzmkc1AES7dYtTywb5nxLhTAAThZnc6VKrpRw1g+eJAz5VATwpUQ+hsdZ9Za2sTlRjyTn+6zz
c4JWcujcmmsFhWtHkSruT8cyGr+RJm/IWLYpkH/5jEWQjPWLp7DeCpvwkVkEDv9lClwyL7kwKFBC
S08+zXaFbENeoAfS+RxIBD7as8hWF5xEtXG0Su03h5Djm62SUgffKI/VG4GwilrY8LAXW/4vb9ra
/gDaNrJjpg21ivfyMedzSFkW76vEOuFT7usIM0ZbGmNojiby1kwrmPyPK2stAEl88XpJFKS8oEfc
xpBg7u135o+RHDadX4SnfpopgBooR5NpzZbYId7GpgfSvrguFjAzFv4bQT+CyJappPtuCO2wgrd3
zC8E2LMAupyoEa2yFVPJIIL+EL/IXIpmWPUz0o5lHvkGxISxTtAkNDYvbGtYDGdQg3DpDGTySLCj
ELy0tEfak6Jo22kEd78lLePUqi6wJaDP8wXehrWjnK8KAgCXwImq2HCDhFz6/IZARF7vNNxZnuRH
R0kdI/nXP2Luvq8jAoi28Ma0uA/Wh6i65LLUJcrsETnwLL81RVwunI7KXPr92bXvX4iJnpJTaIUo
MqeOjoa7t7VsrOI80tYMfVW9fgZQqnEGBKyUZGyV0syUACJOY532efb+D6uQ9H8b/NaVZLMLnUAy
vDwJDm3CJTMHN1Lt76R/T4ZouN7n6mQvct52KWVsQA74c1Re39MY0O648rhy4p6fE4FnNiq2fB/2
B1L5tQLwz3iJ0j75rMouxWSpYr8LC9QWWzy2FmpkL3ccTg21Gdh+CJ7Pi6PhQy7vHwGnOf0oFTmt
Hpl3Si+1B2RP7g+JV+lJHcwM91i5Ac5+KiP08pjUam+c7tiKPSUdm03peZnK67LlhJnCVxQCJRmH
GHIxG2D1K+QDmlDKDDn4DuTmL4/BPTpE/9Z/vr6pqWNA/Tb+aTIBnirkfk+b4QixlLopDSsdUOJt
eluYlud//U4SodzPr5Qltpl6Uk7SnueOYorRDKbCv2fXlZPZTCuFo82klZGTH9l56XY2c8VUbliP
GDJZt7AAYU9YMiEToE5/GLfCflV/7g8ltzrJgZC0gtAMt3nHX41+4KU65a/Sjwk7u9WrEZMSXEng
znUEXRuCqG1BVmdPcMpHLixFbW5O019bKRtWHMeCzUBYVsb0YD9b7P9tk3R54cysKBIwUEMPZ0cN
3iTz42avGs1Mmyl4oKEx/H162+lnzfZbsHn9TcrnzQc2gC/xA8nLrO12nzRMc3T2Dlsd1qllb9eH
mIg0EdKk75dbD6p+CcV0kKZkwFTuai6J1S+tgO3MwEg/ZRmV9WM7J7kjS1E4sYsnf+h04L6YSdBY
rRbcKFK2i3B+C442RUOdjjPXy3T1jlxRUxJ+NxL1r0Phn2IkRSEC9R85vRJJpCwAwUoRL+OBRj92
g8BZ+u93G0WZWd+DaUKFY67DGu/KuyPXvlff9pg6gULzuKOU5WsbZkxqVGjwjuxYi5p51EXt2PAm
NVygWyeSqyZ+HJS2yfBLtwp1kVjBNC2vcNsOW3MClNnf9egtPkpto+t8Z36xolCC0ERVFWTTGRu7
y9dCHhYVsHZsSte4LRX9D0mT40vXRoudjWhQUskHr70ebeI9koPtsDCKgbH9BB3vX5aESKJMQmcc
tlcpXFXO2nTbssdagCGUwBUxwXS+RGONK+Sf9ORPNnaZ+OGGx3wjPgbRKHmE4r229Fhni7jshV+z
hUQbPwF9Rw1QSLeRkDNx1MMK+2o8Juuicq68QP0uyS/YASE9MlayqhwDkKJm8c6Fo1wPkL7NhOgv
0sjKu5Fsd73wCHzFVdkPVPA+C0ZacuJgZ/4X37+P13tzxEDEuOHl8ebhkNqbyW3mS4Q5SmFbe/vz
3wv21lkD7u+F0piue9prxnuUfeSuQ5hZ0OCxiShz5xiTDWLyYsp79zt/eXFzNLkYPG2BOahANuC2
veN4i4gJa2g/04brPPtkSJweY2ayyIqoWhp5qlp46jo4lFp+PoXfdQzl0VSwRaKXKHpoLvwhI0LK
9FmYj5lKNkxPDdw56nOHRLDIYylQvyxMVTvMRpCLKSjjXT4tQI1c7jiIlx7/dS8mVe78GBvkBcxv
H71wBrcu3XeXWVnEmE+CgR1QtQHgJuFnkQ4i+iOx61QPu6RxgvREhgyvZmv+aQ5rhkAVn3YDl0or
8yDeELVhy9pOFNQFiGbx1xN27gljmNLbJWKR+6c2TnM0w+4c1gwKPvGEUq8TYuJx6DFCqKcA3BAX
7EaVW+9sA7Bb+PXUSOjVKgdf+Fy/i4BwJ5mBxfY/V9sZLr42nzSQFOwX9L9T8kz+dvQFFpLr2FcL
kdVWy2oQyUxJzZGwcA+yPKXIScOU25cgO4fn5SqgZ8zZKRFPOwe4LvJjKco7uPzOlm8yLbKlSpTb
1BKipjTqn7DYOdomDCoSCJlE953cI3wvKjTyOgUa9/TpPSdKJgpEwuq8vXNxWgtudQAlpDRUQE+t
8yLpoSQ4304kxe/vDDm1l42UXE6NsTw4UshOtYtBRnVfiXK4Gw+rukt/DFth6hdChoE5lUVGa1mf
y6D7jiLdChaBPO3+tjTcKeCyqZXOc27Eqqz3CDUZogXP3MH/DwhHxjApIX8Ko/sNQxhQvrE1+Sze
Kg8dz7sjq3ezJTJj9sWBYEtGl2z11DdeUDFjVdDrrFWTfkH47Rt2w9UN5FvhYlakmg4kZtWyh//W
uo8tE//IZxckKWeIa+qUDbgiKEUEQoDV5zkwfY+3rybvHzSdrOtbw2+56bkUlH/nZyTKqTPWngTh
hnicSndzQnHKziXWaqLp5TAYKJOmkzU1+IS3TNPLjxN15LQ+XAZe2Llxia/cih0RF1WqRbYmJm00
IFS2nZUczbKisCG1H3P0T4mVuVaNUcdTrr37XNkxdGWrblc3zo8owqQu8SLqOkimGxZnSPKEzM6/
RanDBJH5pIPIObhgjHltI24gcRBpUmkPyccDfKVsCYhmaV1wK0M/mAnFxWIgjxxRULoqCZTdOemq
qPMBaB2NZXbXrxB/yzi/QFXuvI4S7vhmQKjLY+0sZKWIguJ4aywnLu3izaVwu4VLRQosVUevCRDE
4eH6T7axe2Oc/oTNEss4pyKl9xZZUkxcFjJ2DSisMV2N4EtcgBtrnBVBC2HgnQMJc/DF9UHU2MrD
qX3tsxJilaCTAnjlQeGYYxXFmPrM6m8tkvmfe94uU/RlfRs7EjTg9RxGtlH9dtmBv2LaCRVwHN0d
0CsToEAr+QgVNX5n02QsF3t+YYx8nCyKNEdfNMjnfCCQSWBUHNFk+qoFcSwr4gjlsDDhb9dBVl2m
9FXv0lbTzU73VSbL3v9ZFx5SjgXv8+i3VNvLF4HwgrLi8PBE89EZqPpoGw05/T1r1G1Wgwrhbc9a
MXKqh8wOCgdDuQIgoWFvxvo8t2cCGHwXqpEuo8Bda4VwmroakYukuT7CzmZ+r6KBk1YZzwZsWgrn
0RKJPv6/EOZ5Gz+1lVR7/W1CQ48XBfuyNKWpo0iZp4yEQ9I09LFdv7fA6ct+pgqS1P84kNMkLArf
X+9a0iS9PMqCMIxU/5uHjiiTNL7wyvF3kHD+mgSBYLIbJvdYgOo96opbgNuzelsNTWkDOTAijh/n
yoBXCSNeJ3VgiKwNLBi8A01atKdkJqUMED2Kv2DTniyTpQglVtYsKskutzX/mfhCg2pFGlQWHzj8
BpX3sO4NrhQdIqAaM8BPu2XBTubf9urmgHpuYT/8X5G8R9C3xNuKKGtack594nG/o++UE4KKEcUs
hX4+9HCG9VGf/gff7lsCrpFweaBCjXcbyc2tmvHXVRzZn41/4CnUSyJ9Tx2bV3awD2d4W8Kd8yih
30RvZ7tFNyMfmsOvQ5g1VYDqBHZkjRp+71HE1EcsZVoQrYq1TmgMeLOzdtdVm5axRc1m7t8XhoAE
V0YkOJ5TQNfRY3ejllhB5kenGBPP+xxf7YusxeLlCnC03glwO2T21ReYbQo3HO6Y46k6N7Bu2m6I
L9zVe05EZ4r0vI5MDNPAI5D0zV2VfwgFmNZxgmiisogFMRsP9BCjvuIN5P50hZ7xZ19yigPZjEDu
swY5CDr4RotQ2He69iuG7AFfgtWyU97Hqwhbe99HgsSwRDZY2Ztl5c6mC676LP6PyGdEFcYzFDIN
fJqFskyMwiOOwbKVc8iV2iP2v9EAv01SSOYPWI2lvoXhYpt90g+pSFTba7ZE19c3XyCcEfKdqO//
PGlwaHo3e03PgVGMCuwjM+7b84eE/eI6x1ps+VuwLV1y+mbTvuJgnEcC2evUZRmEDKghkKd3ozl8
bkleTc+CCt+OjUOaOj+i0ZI6LCUd+6jB125WJfUFof/nN1AFr50hDs39xvwSquIMzihNQ2emJTdv
iuEDl2AplZxAcfY+B1uKmwkQQVrUo+l+edT93W/Qu5VVDjuT0WXbJDK/M5PBcfCqlw4n7pSYt9cE
tn/2zJb6JOK/8Dk2bxtdedzgXOeh5pskT/kRoSj1G50l4KR5e78H+a0GlRvhBVsuM/lxGnR2T4oL
ZdietDdWOyLPnCtpATCcGv4BZwFg0itLa7FcyJpLB6Ya4oNFN/8dnFUCwvyN7qv/xv0zIUnOhZNU
N293OPf3HGDHLeJ020adVmpfX8nSUu8yMUTp5BFeSIfTwFSbmEs0zQa2g54/Ui/4b/sCMZybsQ5v
foNcE9VykJobihN0YxHrLO8HasajMTVPPsssSrm0Aqd9JYdXfPaHXb+CNvhu3DrlcXGtdVV6yMSl
MoHE68jGPa+E0vvoAABxKX2AThm14ULQTWlR1TVV1iBlK8jr7DWFbDYybhmWrAmF+FPgSV279SUT
wtDzg4yfFurFgzikWtcKZsOdyfDjRaC24RjmQo2xlF314bNQBqU9hRkrD9epTeOwkCJCxj0sRRuw
wKYpPb6A+R3/vhl/6ecOHuvM0JA7LvdkkrLuO+dRHzcktPbEG2Lamj1mmaKOMHmbG8ZZAhg5VwYj
Hs5SW4fouDqdh7tiGPMNMs5FiPRyh/G7TDH9m1oirXWti+NHO+VkcfrU3A74SvfZEY+UAnbpmphW
V/J5pmh2owKdubblbgdhEOcw1wK+sLSrEiE0tI90z5nvcfPg7ZqXEi9i6q0d69Z0140QfAhhgvup
psUo7apbXz7q1nAfftjivbB0wTeKpi9NCUbwr1FJG+V43IOoEkYGhXx7+xwiUu+P5ePBhVj3Sd7t
JQsjmVr41RnZ1Z5UUU0rQeETOVHhk2oYbx6zDPeXgmHtdbc88VEOOgqJomS0CATcITcxXpjW9xUe
9VQgHTy/jcCQJLSuWAHYQHOFgfGMyuAREozOC2VKS+j92In2hQolxTZ2PMjWfdeClMhF2FiyawZ/
rYjzc57uVGyFAGz/a3QAqQEZ2C6FUqwRI7SiHD54Ur9JVIpocswiO/LpzNtVCQOE3/JzCiM1uvRG
ipsCA+xGzUXK5OqtzxVmCPdqVca0hOma4jqx2pJXD/x04hV1E5L8Pui2lSKpnLh5upRasiOC+8TV
Rq8FWfGxPPu8d3tB9JWveJ7PNzbIHKhEwEXrv1qgsrcp+ua38Z4C2PFKKpX3dlp+kwAlXhv5HGQA
d5ObMACodndtYOsOABYaGI4pVdzppTN8FXLSd7uOikfsbVRTQqp+eqcdQpqBWam75ib46EnTR8wP
GRv/kbSFAc0N3cIKLWtG++8z6aQ/jpM337x/HmS66Qrj4DVw240BhCtqzzEmRCPOSHco9otG36KF
YVne0rw3+GSkTZaPKFAQS3nJY2MFYSsewmMBP85gFiUZ9ilS4A2wnfQxqzDgaO8IR1+47ihSJQCW
5DuBRL9r45DC8fNSORrlOi3v8IgmXco58dS+v45/H1wt7nDm3k3+DlkglLmhtcUDpymB3/BFUJyi
ym3yq5OjabfuT6mhd3otDZp3HSj/7qeBzVmQesX+ynZyFulBncmGyf5NpZrS7Jhm3Y+qUaMj3idM
fMMUZMxc7KUDkPEojeNZROn8aIYj3JIhOSLWw0zR3kR1xa4YhSa91AwBKtNJjT0G1yfHKnHb3mrL
G7UADZPjge9ac3ozQ3tQD3Ds+IWhnTWAq3Z4K+fkSDpHAR1ZQSDmtAcvKJ9Hjktxh6onWA1BnysL
q3NT5EFACLYdFy53eWLkq4oU8Ns3QpWvJFphEyp2TwMLmU4Pq/8koLzn6EjoSZ4/rqk9kjobq+tn
KRIZpXFomN2kCR7sC75YK9IxmxZkc32OBRvL3Z0NqeLTgyIEBvU5kOWfaetYxz3SLwCBbfWl/KZq
2RDu1XiASOQyuZ1yt0p2HDQNw7tftej68lgTnDmensHeZuZXTQiFoTii7IhrasMmlLPs2xm5CS8o
Lb8xq/Ny376gXfkeVWvVqp4/48Innbx90LDmsLwAXP47wPXMkbdP8X6/ebNWJPwb3dPj/uO/abDR
uuI2hzbd4/Z5Kcziv+BAtunfl/LUlFDDJq5vXzm3bQdbeJHuXLObkStR64JZXIDkOg+dfKf0Jiap
h5K4pLacxcbVNetG6uIRY6GEe3Fv4N2KWEhCKK3yhHunTI50E5LUeumqLloyYxCThejjtGIcqNcQ
jxx0lXcswWHWWO9SuT+b5lt46ttt2ZDxiUtsDtdKEZsggKCvxCjCDoaITlSEWDVFzqSsgCRSt6Z2
tVL8dI+laRQ3JM4nMklE/W+OobNRUIqcEw0T1RriKumaoLvYG04XRMtJHMxiXs3NOiLrBWu83Eab
e6FQPVcNA0kfWHx1VG3jdFeG8BJMgORfzTh5tm1/BWSoIZKitZD3mVqgYLUjEvvq7WA5esbPtOKY
MeNeJ2zjE+u86vCHIow9PurqQludey8CSM2felofkACGxaoF+kKQRv3A9vAxkNseU7UbWHBPcSBc
DjB9Lg4erUP5Q9wf1W3cliJJl1PDcpqwZUQozRL+oFvEBtxiFZGSANj+O6sCzSqUv2nBxLRcgdqp
1DbKi3hS3Z9C7kgQcrHuOIA3zZmKz2o1vlvwitR7v7P9MdblZhWeyueVNe64m03tmdm+8baqp+bD
REfMrdgUqN2jphvidT5UdO+sXmHw15SUI+Bmefgo7Sv67zYyU/UhYIaxB5ojecZt6BT8wfgnfFhG
gXuo6t9+mU8tlpkFQ+1PZtDzRJi3qXNO6LFzOFRCyhSH/riPPR4VU0BROHQOzkNTyjV44Yr6deTe
wNX/zkLV9nV4qqxdZAvXnZBq0NiawZuxBfm8GNOBEvWz+Lzf91J2Axnh/O49966qjCzF0P5OHEfV
fUnR7lSC+UDi8S+hIYWkbsmVsrD2Oi2RbdMnkpLqTRyHl0H8uT383P/hMpY+U2r421wwDf9b6qcb
CJ+sco/B/z3/1yg5R+wezCY8NKQ3D/D7BrEQhiZmdHHqudF+ty9JwKVi12jRPieU3HpdTdRcpluR
wsKHkwNXfZ4i33AoydV635C44mRRJattwCzkjbSYpLDa7b39xilzg1YH+fzBYOMYPPVf263532mH
RW64wdlLKxDyodpW4eSj3FPu+PEtGqQmR/wr8AQ8Fl4RbbK2yZcej8TmEA7Va/MQa1hxsjDaW9qm
0FvheBAbku/YCu+f3PXXPK2axaTmLizNMj9ygfOfVm2s2Cetmef5N1nsQ22bkl+Ra5jJJA62qso3
4X5fj8o2Nw5YobYveeLEO+8m7rggz4yTFNIPE75dVVhl89Ji9p43n7xyfzJ4NABc4aEUygOL4PjV
RdM3rHUaTua24/ZpDvuGzUgl1v1/fMp/Ld4CSbkcpx+tBFHWL2vLMad3DJFEtsn42JWPe4k5FT9i
dsqg4J/hv2ZRTBpKIAK4GshPEymZVRgbr9HWKb9NNf8Is3kjfiQF8L/5TKTbOsRfGqbTussXzmRL
/dYjGIpFMYimFkh0gw1NvNyeAVxc0WQImoJs5Yjs+3V6tlvQAYgyhrxrY/edif9qFYCXdD9H6oiN
45CYLLY0uss0jGx7io9jget++1XfRlbHZHwAZrcIkCSd3xhRVezkIW189A5m1A1k6PFB8nLjWPm2
6aCjpcSXEEcXDnxZuo0MRyE9oomtnP1sv5v2HnJaWCU0sJhtycJOHh3132YL4N8SBrIXhAiTHBac
XYARFn0Ry7BK9kyUCQymiWTuMwcOlZ1WLmRTKU5CFm32zUgH/9WhmmuT73Ad1AvYNnJSr2YKoH9t
zfrHgD6skx3+/Bk0uoR5TaxSuJNeVG6NNVa6qOVQsUzgoW5a/X+dMe9bMk2jQXYAaVdla2P4sWbs
xRu15ztJekPoszJPDGTx+oAceJ9TfGXr28f72PjIOVqIv99UqpZsSfQK4b0e87nHAesdpHmaQiK/
62lkGMXV6eXBGRz1rnXrTiZZHUNl/cqPxUKFyQCd3J4lIRVTAO0ng2a72K1KuVSrv4grwEVHGV+q
tJgxatLZ4eRKumTfpc7BXgAbZJo1btEPjSAmBDXv+Bmacx58Ah5jcHHoO1N40awElW39ZNTtvtzA
gzqhmjun8Ftru2WZAw80IPXfecBuE+Fmk/vnOmQs5ug5HkjIPeP0RVzloKjlXRC7lcPhRM/r1Yzp
G746vpkI7OdE+7zZinW95qqPhr7ryvarqSbp8NjJXIxng3+GxdLCbp1zb/LK7g46X9VA1plqbTrW
EF+OVo1+siznWHsjaf0iSD/4ZjFpuJa3pDqe1vQi9EfuduFgwW0kj5ltr4BQxxMVhHrVsTJg7S7K
z3s87o37+q8epty7lhvGKVeS4ts8IMy+uRL6kh4ezYL0fa8rHF0ygD/aYoFub3c2qPJwU2H6x61B
9o9zy4Lz+4H3hhuigu6o8hI9BaGoerc4A2qSe99v3Y4L+AUeNnXrsTsfNbM70UyY3k1lBivEWb0G
9JnWUCbYxF3HPdMbpsA0SRebl8ymu9LkWbtGF702sQzNCpbM9DuQW0Q8f4X+ePWeDp+jsuCtTugN
2mWZ94eETNfWGzBQQMEeDAjxkS3U5+Q4uqWJszBbBCe5z+MgBHT8IE54t+HPt/OJPMQ2XwFzeX0l
7/Xd3r6f2ER8243n2Q/7UMW/+TBW/OvZaGgL2rXpfAWGAesl7lhX5jji3onMQrWBxhnycDoXMf7y
P9yn8FVCkYp7KnCQ0leIUT+myAfHb5JPEKBSozk+cePY+538bshtFRg3IAi0StKn07XBJ7w8/88g
K9QVpgfZUaoBCmNjbrcbMK3s0beIi1pJL9LmJ4IQpYgX/Q517301dqRDlfzKIZPhxSjwB656iCxC
lHQPi9DQFvhm2Ama+57Lm4PYXajlOtI2zzOzxCb+OAD/ImdLyg35lVnSbwpNtdzl+i707IvDDbcH
CbFov0KvjLAUqFW4WVApvJznyIHUmHFROe4QYXgtDgBn01ksB/JUqzviWcfZ9o+JvhZc5leebO7H
rSKt78g5T4KLEnkXBA1jUQyMKrj5GaaN0zqPbN7PoKti+y9f13Rf3Lha/hqob1GMPAUgYZNYJS1+
jis16M5kuCYfip8Y4klfQ5bng4BG3ZxXQTGWm1ltQTb7aw1lI7y0RN7666dk1YY+RE5n2MZ5r9RX
NEjol6EjGKeqUG6YY8ZGUn/j+LjhN7XyJLiwftpZZsyOB0Cdr6hKsvdjQrKXqMlNSP0Oi4I3svTF
/w/uWOvMpAR1CXT+Khfjda1wZdsqQoaol4rMb63l+yHQFWSrkGpBA+4ErofVOgP+OlgdnZRJB07n
CNIF3mZlBrEEVYmy4jRtSFX73AjhdPJcOVrktOYfBZ94fyOwoSoVDyHs8HWJ0gjpXR7HYdM/q62c
rWVqDy1VMA3mqFAWeQbEEdI6WQfPSYzZbsbccXQ5ZhIOKYnCUVhXLlm07yIn7PIudirdIywgioNC
XDmfhA3Mo43INNeBRH6X5mAHatlrBxt4x8ui4UBDilpE4JcHN8NR0gmN5D+UbXA32pJZu0mrpqaU
QiO2QfPKGok8jAjDCXk1G4TfZcfPK0TF6jYi6dfPwbEFUYIbz94ccFh+0qMXl0mhGhGz7xJDj11j
qCsQaIOX5h0lTHtscGo9xnosOelJzdMQ7DQ4RzRxxyOBWeUMmntfTLhJLRbu///tJ19HRSpCpCSb
QP/o3o4NlU7xyroAAHf2t9nMbTV73VK1ikjoo+1brx0BeO6SSQR8onXTS2zzawsbDsyn2ee3D3Om
/kUjAT2g+vdWj/wBpo3Xb9sOwtjuO1tIxFmjgug/wx7K4UwFlPF9EthHLddwA97Qax20Rby9jNjx
X+9yhr4guPoYHkchj0neeUYrMiM5pAJulILf642pGplu/3jTxm0fSbqrKmQY1kVhTtcal9ogn6jT
5TV9CtD+n5w+TATkAmjDvDNuKYrBdaa4yUyd/fedx1F/7fLV+eFjI2nxwmdsehp0kLPjLY69hEbr
xtAmsZSMg+uQ9YVb92R9iH9H7TQKJblXHkdFC7PikyceIyx4Dq8/XdfLs9t7YsEqyO9l/kZIZpIU
icH5e02n7NisGgWJqe12S/1/80mHc8788WYnPcnNNAMbbHcqZCnsOtkA+kTw0Z7A3VxZoS3le4DD
TrBIABMah1ikvsjHXBUdt40iBq3d4qJQjj0dSh4zIYi+iESrV0sVhwjRR5VaEdkET26JyBEzpT7W
N84crMIFMi0A497kUCakmL2EEn2M/pVfqoBYeAtylN5QtfTwUMve5dMiRKMqfmtjJuNgIbZphUFG
IYBWnvmQt7u3+WfAaQ3vbgio72uCLS4K+HAQoX8Rn24sUw7D/yzK20184NyjNtvWBjku32aBmbae
x5Au/TxstSkOlWVkMOawgaB/mfpfAaHqtVLnDGo8deJ2Hj2I9ftIAjC4TqkdcqnWVI6J7pkSS4rF
zBkCffLPSWrMt/PHiIa0yp6xEw5bJ2InE6607U3/GBfXwaAMrnxFQk8pf3MGZ2aZ3WS2hS4zpXnm
UmaHE+ZIm/+rYe246kc0QGymwXdltnrdt/FytW3a24RXsj8m/AegmO2enP+7v5N9sWKMslOFoBEX
NfMGZXlW0Tt/b47A1TJDIKdKZIN4yvwR/uBSrz7N1SeOyClThYUzne/E7TnGU/BzpYsMqr+RpUu7
NtLLKUHLjBFZZkwGtFkNtftEZP1BQLyOFujh5/1sPMpxezhJG86eiaOoFP7e0cgoHlgCx2MUCNrj
6Tz5xglNjz+wfm5ErZvXrakg5RCGU+7lSrcA+md7aLZL5HSkgGkEfR4qxdkSh8VA8VLxEUlXVB+j
v6tV7tBXgd9dKmBo24kK6TXqU/n3sIzhwbsraaZ4Ae2QHXoLR0sr4iL33W/+PL1GkokYC33QgcKl
/8b9Cc8O1D1y1k37Wy+6l2qFmKgoCCIYnU9kMwobew3Q51rbKDST3kqWFhOUZeucCOAsOWysTgUU
Y3LfvQFM/sAVYotZTXK18A95IJeYlYXe7DhiTdkLsm+7OmlYHczbbAqAJTkhXouEkkRnyiaGumT4
PTneemontFxhPGsDI4V4lM+2s2p5b/e2OjxYBSTUeUdKKRCv2rByFWANHF19iY9hl8YLUW+k7ePo
x5xDsCKDtFueR7vVBHwGYcEGwLzy9ML6nbSW763JGunDJ9zsm3k063qy5v1SABzQDE3xonJ2Gavs
mpXlknFBvsN1h/1dISdG1rsQvZS+eONMpjBeAzvJsDeCR5HINdD67d0Stbe8Y13giOXxISx4xXs+
vErktIRQtft+qY001OFyVlY2c5e8VrLJl8YeXORh/QKSgj9OiQDhhvM/C0yHK5ICDa4Vi20evQdg
w5ot8PwzzPEUwSDyjlK/GVaTc9TnOWu+In92BEXOLCT5aH9iunaU2o02nHhxwDRfwCQDTlDcnBCO
9y74F22OO+JWrtiH0eJSPcFT5YsEbfJ1DgVH8d/6BlFVMA1JA9nSWwEJOJ1mOBxFJnPMtEOTkTaJ
5pqKbqUFTojitst6K1Rtf99xzaX57xfkDZU5Ecw8d8Gk3k6NAiXB05e1ohmGozg+Ic/f8hTddeyM
7uNQdoFvoPptCkVNKeN7GeUKKQI6BTEJdTflwcrUtDvLncWlUZiCsoZsFna1YTwvpNmKcZfPLS2t
hqXf6PPoukE4X3cI8JhgajoLnqy0JvmtQ4e8qiZBn+NHi9WrVAMzziLhJRPJwzl2Ba4DZq8AIV/q
b8Z/0TQqFQO/fe/G+hidmYrFIntb7mzFLIJqnPHFPf5fh4A20up43wU/9jUsGM8FpnOo70dDw5A1
Iq75nkQq595jD8ClIoGAy9XfHbugGIlUpLM1HfKJ1u4alzBaYiMEzjhiajwvkUGJl1sR7ZhoJ2NL
vMo91tELvY4P5MlwW03zRYzRsaTX7e1LUvhrJCfniwvLaPW5eLvSSuzMSVsak2EC/C6FbnALgFky
PyAuG8B6Tq3D5T/1gzbJuEriiZArGLTFPID0DJ4d/GRwkqiqq1JARHFllWfjTzrquEce4QVOdVjk
IkkFEU5hrwZKcAfxd4RZzNug4wptYMx8HvEDjnqhhyU6sL9+2SEbQk3ViAVWpY19jJ+zWjydg8VL
ZR7De+oyfJoRI3wrM6pl2l7mtSIDSXoFVLs2/2c9tcXUelRiFMRpALKZWTOoghay+SQufVCImhd0
wwH25PXmfq7YmtGdRez/eJm6Nz/BEkP/eUXxR+EKP6S78/x1xu/F6L1BX2Fo97t44Oz1h9eXV1s3
DZulr0hhboKcpnKIlH77Cb9if2brVEoGKsCGffB23aqVejMbiDpIT+ymJHtoJ8fPz2m4knqlTumL
mmO09vMRR4Ux3j2quFTwYBnQP/Vv+XdLI4eil53nydsKoVlriRDFp6VOEd77YRUk76L5G6FPgT8b
c++kZ5XRsjmorKEjRLtheNtpO09c74o0AwwXu6XGwC7plA8cg474I+epHHOHFshDSPryhzU0O9qL
lEny6wT5kcNnWJeiv+9eZWqvAMZH9qcnMEAj10qvlUi2VlBN9RjZvADbRE5N3AkBB93y8q40QWGA
1c9DkTJ0L4zEspLyzid5ks9rGZ5vbQ/btwhO9vz3aP0bbetLzJ/PKHP3Uhiqg/RPXkkmCzgC7Lzg
MPYKIMWFgq7IZfWiqwHqUr75NVcTT4BJC2vjB15D4vkyV3k3CcTRb/cp9/NhoG+wBGVUvVi/zAqM
VJ1owR0FvpAmpfbgyxDzRHIBgML/C1NeDn0Ze66t0k/dOEqY0cqCE5CYcvU1/CMUZRJFYLxjF0U1
QMrrqaIQL1c+nnSvSOoVwctisRWYVsA9e5MnBcRmkedvoZFIH2fO8k83w/paC5iD4diCBFjN8Fd2
MK1zs43cTA+Cm3moCzlMxgRrv8JrVY6FIGKvLqC0bnzVSK+xvKu8ozJwbk2DXUTDTQp+Gc1zpvYN
HN0A1exoKe5gY5hKu4l048blWmtI+O38Sf/BlJ5pur8Q0U2ZtTHgoG8HhfbFjLQch6pBYPvR/iI/
ZYxtsIUfIpbvdzIsQttANl2/Wqu3N7iLHLlg0X6JQIXyc4vr7bSRG9IowZ76l02KAQ317+0iGApK
2wVJ+69bhWLpk9PXayFTva+yEGn9LfnURdBDkIY4SYqWTBonJem7CbOZ1tbMwAC5mQ/oXhEBYf7x
/UTTGC41BZWnb1ZLPcQ/A5eOgoGhXVYZNhKFUKbecrXHeubbc7cmsT3uzjReNpgaUoFwkoC2pSRU
/7YSDHylYlnLWvUGsJemIhZj8m13IQ9jIpnrnHmZXUo3mAgM7OiZlxlPNVQULNzzq3ZKcTfUN2PW
QIgERhTjI78w2qbD+PxaFtuyfkHNisoXSR57TsLZQ4xv6WbWz+GxpUuQWNUqO3EbB1Oa3voY4hkW
DjT6YP+lgUbfDQc6yJrWaNrFG1NK1o2GKI94EFNSrv0b9NpXB4Xd66rJ34C+Bmo41Jl28lGuc5b5
f5lkXriY9N9iyibUCsuYfZH4XomR2giffYQY6p6G46mCWzbedlgg6VLWSVUF/f9EwLaDRMRImadg
Pry1oLaG+xfuU5LZhBmtbpCzAKIn37T15F48FA89AhBfAza5S8Xw4RUEnBtUIPrjDMNmknOqnFyd
uAreD48T/fXpPOeXsM72zijw7tHlqrak7SrIVQ/YY4R0nhypRRBkEuowHey75Y78Y9G+RSpstDPE
bgPb05ZDCSITlPkm82Qwfxj1DPc9DfWeYbM5vfPuPyjnlzfNZ/3HHuDBwmXeSM2w3ikWFg2yf+z3
tpFKL4d9q/4+k7xX92/18hLEt+330SPj1Pth2ljZulOYvg5W/1nQuZK8NoIgQwqo76SDa3KzQxEY
8ifQO4Ew0wGrQMijwfCMTKszxhlqJxNazOYpoQNrDBDMvJOd5px2IEP81hjrS7EYm61DZ1zM8Eh6
B51ZOwcY0/eFhY17FHWgatH8742WQw3Gi6rYArQDLFvluPTHvBRqOm1YEMU1IIB0ByPcYp3JLEfx
vAmb+M2tt8f2ajaM/lBFvtPk3a/B3MYdDQKBaxnIvn2rG1g7lrP+n0LeEXjsAx1xLiQhhhUEWvrf
dEcXJedYjkgLui2UyTEMhV6ZsujRKiiazrOmqKT8N8KSGcpzS9WGsn+VSRNrnqzvmpUiRwuzHYI6
773wfIeK+/XQC3/fGlfvL7O0P2Tf8/b0ooWq+IMEJBPhwmUUD6In/NkIdwiJIVBdS5l+1x9NT16y
mwsyg5fBBK16PdBdQWznhqpjBxpKTfptlN+hI0dmpyS8X9j5ygtwCjGQNihhuLXlswLfd3+H1zPR
Aqirb5e80xSiiu1L67DBw9JEKfpwjOGzgbZZ6HiilkvnFvAtpqrYor1hANeJAqx91bevljo6gDuj
LP9DMFWERn6WSBWgatRrFG9uaixThnIUaltO5By2u7uZx3emT35ubs7N4i16T/ZMhYXXZLScqYNK
wE/Py/clmUiKNdK7O8E9UhvYoFDLqqnfApleDF98U2ZWXAYHlKMOWCzcB6rdr93aSXPt/nCM5dG6
ABG8nhyb9vlJnnfPOAECOW+Fd88q+k/Xljm/Dkk/sNYluCXNbjSm/WEHkJIZDHlueXLs5X57LkFT
3TOisUskLHEoDEnHfkwNX+I+/nBx7fYakek/CU/58wnK9RfvhAOgsBjX5UN2fBLIjftzkLkjTj5w
27zwHAmCykpYxf2fVEvx3K8bScXWmEPSehs1NJjxLkgWzswEGpnYK2f01nmhCwv7bMn5DLwW4DnW
mqgI6bYMoneSnPAUoTVdrk//gpf/QErwaQ8AVN4wwulZwqU7K3r7354TMpPjdSSyAGXsReDGjmUF
TtoVsYI+bRw6rY53wpov368Pct5vuHKXYUsfrsksNRdlnxdsNUIqv1uDSNaeLv9YaEt2nK229XJ8
yujChwRZEa7RF3FjV26t7+vXVyDB08N19Wyjwc2aCDtzbAv1FTXug7Gen7UQM0r+2fPFvm3qiOyh
jqcqbjnT04NHvjFMLV3+SdTWJEwywLyh2tZbDxVxaQuob5NCNEVQSXBpoTZZQDCumaZMF72Tv27+
ZPGrnYkTCHoLGg0Yj549b5pQ7M+DNXePiabCtUM/W50x2gBfEFGVOWf9nMCH1qFUJLHInXPV6YQZ
EPhrR0inksiDpdHtgpFP+MwpWpg0fSKLQOt3CqfwzaeSV6f8YiW+b/O+inMebAAgKZnbcZnT2qHa
7lFJFyrSLBDqQ3hchZmS0SqWZijJK1Rd2X3pB4mtdbkT0S2VzhXznZv9qzCnhzAGcnJF652Wl5ia
X6x7P+UqcxNH2TMwE/0jmvqMocYM9N3M/d/O5B8tDSGO64DEwkNxnOFo1axlZwpGBFCK3PjGpVBz
oF8Y8/My2XrjVZqrK8FeqW2BHCc5vJhNKsG3EXf4ydtAVP+Pk5bS42JQL8f0VpMs6BEDLgviLDDw
XAzwagxAN5vS+p7p7r8KnY817zAawCL03rQnx3WLxnYXqIwL5dZJTgb6Oh9JGM0h2aiT12mBoMwo
gM1/ztJZOXrTCf+0MjYcSp7FrbcQHgU44hHXZBcBRXWTk0Hs/x8sQs/8g0RdDskQc6S5ey7bd8I0
4JnaBqFnuHZe0Ov8egi2sKBCZigyA7ax8puOp6KLjLIjPa2Oh7S3ZWWqM5Gz7B2J9+b+gwpU+crD
kzqLyYBjvU3wQMWCnCcpeguZ7RpwJRmfreuufk/kYLpNZ4GPcgkRzE90o7kGTCVulWLDu40RmfkI
LwvLktgm6wUMG9binsWM3elcVA9+JioDbK1G1U0PgUdn1UcmCv7PDRbGJkPfP19YREDtWWfUlula
cBKjAxB+J50r561ar85g5iD5HlD2hceEcl+YCIrsy3W8GKUTdoxD/js2kERSxgtIkJV/YJNaSDTK
QC2nfZpu1QtXk7HO/YqXz2TO/jCZCq0a4FApcBWG1AQhY03ldfCubjcixNoY49SZwkUsLW3oR/o9
YPmBIphP0NWRmJGwemUCfvIVNcU8Tn4CoolqGN8W9LEM2w1og0FE5Ha8GHBWH8e/jvfZ0PYfp91G
cyZ37qpPviSzKB3RRSJW8x+UoeLxinnYVhclDSmdFddfj94FTxcCA1SFkvk/H4ijJ1l/gwr/vcQN
S6QM9MrKRLxB3mYtzxr0NX1IHt7UfgwYi77ULAq2FktBpDJE8rf6wijO/F/60otyhk7/ZKxUnKPw
Nt5g+PYf8DPAzdZJwX95Ru2qwiX9/VKB2na0dgncO6Nd+L5Vq9mJJATlySNh3UQO/fg6fqt9fqLg
aicMp0I+4n/TjyHwGrxIKg8l/5xgfuBRMKOWeR81fdq4NCCLOS/k3H+AqawFBmO3bfF0XwwHWZlv
m1D6nuBlQ7h6cNyNB70E643Mtw7rst1Sc3auClQGzaWxFxagDw39BNu7AO79pmhSTXaYaUFztOdx
w6wi0VA/HY2monfLDHnx/I3Fuo8gsUIxu1ZMjMnqid0r/nFl8UK5sl+GCRShyb+IGQrw9eE/rd7T
amK6x+k3JFkjPYtWptaEPz3xLN299Xn90qhSprF8hlR2KG75OM4cZ4Ax6VlEg8jvCNkfPntvzsmV
nygFtcOYNLbU8FDdifth47quEdU3aMsQSk99lNGEYI64GsEylxos5A5MewFTjHahClstvfKZqT5w
zC33bQJWtCz2y30DQIJm9+7mRbjlMuaRpMmY8HxMXCkWdev1UUpK/boXkeb3QFyyO0hopIv+gTNR
r54/NnJA/dn8eXtaUm3YFJLtgSIOgVKLM2YeAInk522reA8cUm7OvKGHRxeg1AB+w7d3tOrkF9aK
9oqADvj9raeL5I8rX50vwPrUXVRkZOBheB+cb7zgfo8YRBTGWXZEjOCCCr7Xy0SXZ77PwsxGCgpp
FbOsLwMCAzMP1XMzcastVV2as4CS6OMstcvaMfURvTKpVbAbD+SNS9SO2Yx2CeqVMmhonOt5Efxe
b1U12AEfIS+nkADON/w5FVd405RD+iChPyXiLMCSWqAUvwzx60GMpu61F6fSy3zfPl/mZjKHGP7O
aQvEsgB1apw46AI5j08k2c57SiLsR4avbw34L8wtXtsVvqhN2SP526W/6uT4u6q/Se5KGs0IO8Pe
Hqfi61hjP07VNMOacSikM6ehLogbFq8OjcGVfWyHTbMhCNO3b0SBWCRK06pKNg1SRapBlOcvBE4G
zVRyWt+JLXWFNWRTJBvc9sIVy0oHKrpSSYMWxBQdVmns1p3c9KyWep793VU/4c2Z2NlGq+GCUI43
JONuxjqXtZgR8lJnUMSVv9s5zgM0oaWMGpPt2X8PtAtoqUd3+zmpC+3KdSFJUYdpyVxvAwpvfJtI
81kw7JwYntQQLV4J8Xk+X2o0QBE3sdnUhN4mI5/+6lvgPkMA2QG+CwZ6oVYejmKCjcU0/Ygav73A
xhiJXXSBbVHCpt8xoW+oCXwWk6uWunNqM4b9bCPXK/9JyPbRrhTkbrX0MLlSS9zSQy/ePEPZSF3d
y8XP8RmeIRzv7F6GlH7ymLb2OmJphL6qAN8+C9T6CDFxAppHXOMCKkJivXuLab79tjquK1KMJqpY
JFJR1T28w8NaV0GghnI6i5VksfdjZZpQE2EJUyTKq9SXjvCr+83wpc5nsOry4hC5WM87lUYmcrJp
z2lgCna8qwAZtp2OKCuj9uR9d0/W1VLFacJhN1FYy0CNzZODbg08LM04Pj1RIONQqsRS1Z0PzliO
7cezirHjXejOOEao2ynmpUd3m0slIu4BcWmmoH1EdP+yEzisK5P3nGD9ArV9kb0pVyiUvJKyjRrv
WWyaSbSsWXawTVZFmjgUmJpjceNhoHR8N00j5X3ERDcjQuUf97DcFA/2ziFhld4TP9ABZczdU1ti
hYteh/taiajTheWQpcYwL4/nAmAOphjjKoDVISokiqOBT94JRVB0AWAku0nnFLMTYKw+xU6Lko0M
86KGJZDTB1rO+0ZYwpbB7iLwRWH34wYW+aq3LkTrmP9TKGoVGOFry/1uO2ChAlepkF1FpWnZh9gD
g5IksPcwclTWSRG1r+A/eN0uLqPck58zXrMVhq7HrldCnDlxTGFa6D7QJoNDC2NgJLkNjOm6Fe0r
cxvWjIWMksAIyWSIJxZI52FDQ737mxtyO/pjErL1MQbKwWUMkJ6O3Zkfw61qvpm3tBnSGJo4sdjm
YZP4Y0HKAaxdkrqezOEh89HYBY8Ge2lmCgjt5hBrgZaL1W3d+putEa4UW3Q9eC0t9sTBcvDa5fyb
8t0hI66KN73IfMUX146i3GSr2zvN+4cILEANkVUpgGEdbfo+Z5EZR5z1lXN7uHPN8h7l8SEr2hAE
jF5OeCMl3a6gfBY6UJP8+MhSrjS76AFJPwOcFujgvz6Bn3NAtV6eot9OuOVwE29pcMsLa85av+Xg
vyKHBwKy+W8axEwzSFn+EXJ1rBVWKE+45H0RGRKTETnrWhwHuFoy1OlaiZ+dwYUhclE8CFxPKi0X
S90hGTO60fXBcPnPiujbciDTd9MMlpP6URTA5WXzPYDaXGMiDrvrwFtaf9WJmSbW+clf5nSqtmGx
ByBtdv6KBrThSl/nC2SjkisrC01sJ1gOn73Oue0IHaK0zvtZuiY+iTuHEsPxEEQTs4TkAWkpCZpW
JcP2omluCue2OPew+ozIRqxTcGexhiFSsBqiVboj7hRHgUCqN8C8FLrMFzkmk2vH2PjvG1c8nJdc
doDgS6MufX11vUIDcYVjr3d1kDctG6TblpiMOAFH+oo61+Ls1Tvs5CkisyfjbugreRehhxEZUooo
V9kpez54qLY7znQaTrU7Uug24SCkaeNTJPEMgCJ1yP1ezgVsRGbTdeO9Pgr9iAxtO9+4iAA0tW2J
AUwfyypHgznwUq5MmY/5i7wsLHjKSOhS8r9ZyOibzaSqxXi9WhXAucVfzcFI+ScSlAUo8fKihQtG
RMCQITkgR8Je8x/qiJMqkZE9Rg7lqgSidK6ZBtSlO2qa6DFWt9THuBHtprS+GtNWEEegU4nN4KvT
rXjBwdF23ZRVAgiLkkBq50BnOB1UEVdaGM0t95VIFoyxaQPsJQOHW1FKsK0UpXpp/zmGzorRdsHp
qZ89HHXKoomOX40VGakPFzYQE2Rw5/DBGm2cy8tOk6bqvO2mzMsGH+lxEe5FMdZgDWEfwA9PhrCv
IyWMh/89XfcrLfk4oRYa+XZ/RxtOPWSwJZDzETAnAamq/fDbxTIO2+aAWDkBYAh/Pg2G3xMGN8BZ
+HExeKDMbWTjxsW88hfsmUp1jA7fS+8bRvv3y2lH0fJTOEt4yjJRyXgeAGmL/O8m1bcc/96YfN26
3Qfk5hhlXTr0bQ7YeB0XS4xNPZ50K0kFWQJKIMDw/P/6Z31gw9DFdUsqCfqxd7oiNSoSLWIFVepo
fHDIbyPH27OWVajC/wD39NkRORXKdBELjGPO/BKjmMPPs6ViUaHipHJHrv2cEgPyuzIGLlBHnJrc
iUsjIG5MVEBC7cwpxtFMOrpncRldpxUov+Cj3a3HjsxQWgwhZjeMxqO1PV4wHi5vRyaBW8Lfn7zv
dKtlfL6dLK2xsEQbG8VotUGux4qQ+SnEWfW3ZBkpZihFD4hXosTgb9Bdfdcxhq72GbCZP59I1g3f
foNsuNsELJ32VcBue7OnYc4RxzJZcL0UqU1P1xa9x8GpcpKDBw+6elwh5YQt354noBTok6zhmyFL
+610Hy2tbcv5WQ23coXgY0+ToZ9fcpGU1f38WQ9KuwKA/JBp2OeLlH94B5IFV7sN6DSYVrUR1p+J
0fr9A2AX4UoPcS7IkHG/gb8//GEyBVY+f/wmusH9fH+lS/UcFGPtNc30qBevcUHxmiFjJT/+0D1R
ecP6RwdQ+volNwv/Vw/KJY/yeVx+Ylk7ejpKYLmv/StxAOqubZxHp4j7NH9mETGZ5Q5gytocaq2E
qZ0iQYoubvtvVEoTbv2Nl5vQvIezmjd9rgRwROlU6y3jNLDUZeF705Dnv66vZj/G8ZVZuGtaGkoF
h6MoMre+oBR4evO3QDgdbDVpiHqqlgo5joXYl49SGJmMJEhim2yvqQS/9jbT+TvuZaOkCiBliav3
EKI0/cpJqdrmjGUAqC89BCFKMmpkDJ51rQT49RaX1kabwC8jgEoe/WsZA94kYk46EZ+HkLsoHjci
LVG3vf8KaQBIiKelSNb/bercb65IYk2c93NLPFUu+AuE+ZQkTE58q+gjRuEBcDyT6xmCPD6tQXxU
MuB4NdiFScdFrwtw+nzNlZwTuEroW4IjvwSxJBQIN/gPyid6S6TZZ37crUYoMQhoLNEVu9t6nbeL
KPAtFZTkb4cEjZRm0Uw1MeW6CbiP/ThawbUZWL1fIY8WHiIs6vG02SsEW9WvuwaxD8qWpmXLONUO
qd6ZWJGXZ14R5X7M6eBZ785Iw2p8JrYxvpn9weOzY1ZvL1kdyOxySXe6qXlOQ1+6RIi0Q1BmdNXR
y6sSoztOU9iaviUxa0OrfACQPsnzhXJHJg23QGJjmaGtQd9RKYHyb9x4L/n1nF/RbSXFNOj4cYEk
HYiMxs+/SYFCxunYac0hlJB4VlUBjZaBpwdjiwTrBm9XQS9zX1C0YevsUe9iGcf9Knh9XkmC4nZU
N/UCRcFOdHWu9k7S1Zy6TcpOKBGWnnYxnsgoQetpJfO6CpR0pujTmjmhbG88Pc/vF8VdyVyqsAaS
QRcFexyjBv95L07oYDocDEyTCbsagMudjsTcR8M6AuX4wf0WecQLVW5ESNvwrFHrDGG5kwSRxdTP
g7QSHJ1K+x38WEI/u5NDCuLYAjF+/kDD34Vdo+r+bEf2PNsN2HdDP9O+yXoewaktLuWNm9xWbq/5
BZEg8DrbJHmkgZtkPP/WE11GmpoAf+PAXx+6bzbQQbToHrKdNlKmp+qUSGRCGMI/8omf3d2Ulvgs
jJe1Qwtot3Za7knybo/O6d/FrNn/hGwT75npQmOWxLaZaDGNrhYvDYdj6BksaLI/9ajm1Bv/cbCw
nq5rzioTZYaSfH4QmczIQRaYEDIil8YNhYB01tk0p8TXFa23aeWNZCWNnBQuohe4QRmBLmdct3Qp
7vKwqKbzUgV9xk76IqsOlPdAoX4tOEgVhaFyESVcUP1tnMal3aRntvEEA7986l9t4q2NWIOWDiHs
tCl+sy+46AAGx2U1vmICP2tPijJKskSNVU/yBWUzVG1wQMBBO8sF5MTovK7OxGoiPveLeIFOhVHw
S922B+SSrL1zE6M4GwTR7JzNL7Decum36FA89XP6+1mbNbHLiS/IlLjw7gvCmYJS3CP2Y+xm4p7D
TK+gIrKDCsgg8tuyvVVd4nJzH7Jl/jFqmGA5LGJcAv7XcxCaVO3w65W6Ftl6swrJ4krp+Hbdk7xW
X4BKfIlFoorGhbLkKcVWrn8SRtisavcfjqgG+vcTjolv9q9LtIXIrDMbZAa98XOo1jn5yDyYuM6G
+YbN7YqyupsMmmN2bmGhHwr2enyU9WMEZK/8s9UQHX9TcbsWKzsalBKKuIEhcLSxWQ2aYF24Kx+W
kOb+AjmsSPP4wWuYfJ2prX9YfSoY3fcq4mpYW4nBsoQe2COghmrtj3P2DAs7KltHjgWCvOK3nqQp
5h8mFkdXmx7fs1iVLDLG6GUs2ErdNiWtuAJOUZLX8d0Lu42OXAENNI1VsWz4L5lIlvmXpIBCuo0J
r+vjhHQQfNoJPn2jNcXkFD7E/1KM1p4UqBj7YJpYbqZQ7x2TXpBVhCdUqlTylN1/qu+WJ+YpMWeI
n2ua3ZsYr0iBlGfi24UH6tAx0hYotq6m2f/JMO8xKhgK+bDa8AGMq+dC8WTeLRi6Nvkq228b6gaS
5cDVN/DpyTLjSkDIqbWEvJvqYC5dtPm/MyXixp0ZCnJQgTD0D1F2BS1m6rDB2ay+B0UCSUYKmwF9
Y+K9T3mKaDuzgGeC5iX1Z4D1x2IcSyeZxo8orIdGb20oW/Pe0ydEfCAHKRfKQOqYi9s9F1md6eJT
G68dS29Xe/7o88ULMyVz4c2yR4Cy81sIm2W4laW/uU+NqwmZIkIJyxcr8xbtLbOJQp/gZrg/BpQI
6evp6QTppXiy5Hc7PhjKv8xxnnkSVl8aLw8nBIVsDKkmg+wcL+CmkqDAbVZ1wasX1FpKoh+g77Lc
JDeNswunSkZT4y/tsvEvsCmbOVQ1yFQ+5NOtMcz15S6FQBWa9aajAbrC8SmbaSm6GmqpxDHOW+dk
FfXq7m3ufbmyE3zuEqO9HldGUzQJRFewC30vfUzUsh5xM47Se+zWiQGZvfFGyNyk3mGFLpWr/G04
laOVfbBu+5kSLgMSC2+u7ds3SAG/p6kVgw8HMbqXuOHHEuwWBZ7EgSSrUWBwgW61MCSUW23nPTJR
gLm5c1OmszkE9ZbBxarCCj+Yiah8ejnUKUqu+PlUL3E02+gwjpEs6eORUiuktPITJ+ejE/sIPRUj
c/6ZfFOXHKCOcj7h3GuIu7C5QyXoj1NSRGPcAafJYn7OhLTgNR0Fi7cDBwna7MzNU6o4y88QSCIw
bStm5qADOLxXjgHorLyxoYFJoS8ujqXsCWFPS7AkQoI3PakMcI4P4WahNd8HAdIPtTdJTDZzUJ4s
k9wJCSRz8EMYDUnZ33gnIXNi2lXEl2fXeJrNOI/XbqR/Crh5OI02Yut5nFoAGmuglcWxd2oss7iF
xBMBSlMPwfopgDBizVWuRkLbX17cxOuEgYybyqIPXbsFMVbZlblMy18XLBPoEYvr17yy/KOCnND1
dNwQZPduH2qPCFyaJAY145kAk9L3BFTKozKbmNMfHQ6I5XFMbbkrvcgXyhB1YyD+gvQK2IbS80+m
j8V+j/JcWzpA3ZO/nxUexpImL+Dr/b2F5Axhwqx3zaYyX0+Wz/gkog5MHmFz3gAoVxHPBY8fRWVu
C11FP6lYKaeOkKekOn3gmMa4wCDuHjEAWXxb2IgM9owKXaDrTbIWtpcs8AGbgSdyt63Xdye0Enz+
SEGhmVqsqaCqicQSUojzlutJ0ilTRt7worIw3bUZQ7gLRx5mYlE6d017vfUwXUGflroB3hDvvy5e
W9NnQmDHdRRoAm76l4rPYuuLWCccUonyUiIbUyGLumbM5ZPGatuOHBWiGNlq2z9niN76a2fief6h
Y6QNBo/xZtmlYH1SLJi7g84J2Fbj1KHqcE6hd9e/2D7oxC29mxrfAoSnlc6uzlTGCsO0Qi7YHpBZ
bmqerdFwLcgV4JS4D56jm1gevPU0HU5IqTmhEdBJnoDFlIE9UpEaykHWal8pGKJeVi0CAlr6wP1U
p4BnvJLTiZxhgi3bO9bAkR0f9re8M7WUqa8BoVAmCjEIJ087hFlWDE/K3Mfmu/lmY0rj16T5QFGE
c4OzarVBxhh27yqVQ5OGDt+sEwYuH4OWD5j//pjKX0MrYOW/ebUUnjQ9HS/QlCSyStJ8t1BFyYLX
ozYV7vqPrnA/9Fez5SZ5FyibX0bIQ8CHBNJVBsveGXr37ekaD6DM1BbyDvzX2Dd+e8c0LNOEO9Fy
6/2OjQjc5ITWDESrz1O6QFI6Da3HhSpMQnDlyZIwjh3t4C3llHXOriN3UYsgPvPlbo69R9zMeV60
4YHH2Wjbl2uftoG8K1mPx4SIj0PCQj6IMFAXJv/NVtSTgkrmpoP2tfVqcCjW7Nd6WvOoHYe8Uebd
5E4N8yhRmLbsQ1DB6omSTgYf0Kf5iD7Suez3EjJKLnKnA48KaT+WQ1/es+LidPgLaexhcrAyIljl
leuLQFHZyo/PtfxS7stKym6cXvbPyDZ0taiph3oUzznqPZTBHbiwYCkfdsQtqno92YZoRl3o4AhB
B+FXP/QEBNA+xMjv5qUrtaDtATorl+vFIwaK/295oW1fwRDceCyualpds0Yx+Fw/0TWwNoKYh2Vs
3icV+OLzRLHRiyPwTUU2nY1Am5Tl34NSj0xZ67XZumgqNUggbN+ak0JSWEXiYp9Nfvcg+8mWNysJ
ocO9KZAxrSTspWV1YN4jSUl14hZPLaCX0A0EC7AJEh0fgyU51AsWyMOkwiXT65vv1h0gABXBvbZN
JgX43COG4GEUC02C6M/aYOPuKjff/hT7G26CspVGYMOXv+pEDymCbeNHxDBQ2JOewYuC48kvyiRP
AaUXMAq0aHi+FifFSjQ+VJwaMB83PGbVOOh99WUuDsmH+gyEXXr72CdVg9wZSPix8aireo78zIv3
p8/hBexdAv1Rq+PHEBaMIEyepcQ8+zQbz7+HZ+GVmYvulIMYauck8D11kcPzG/cViQXL51Rtt7Jk
lATdtOG4KmR+Pe37yXP1KRYAUGtKpqlxn1alYTiE5Qqy3eKQYNJkbNXjbWqMd9aD0c9xSn5JphV4
fJZfxlRcI9jnoP6AVBB/tjlUMXUvM40v5gBJXtjbrWGOTjAmdEYZQrEAAe0djJoNIQ29AdGKBkyA
yk6dD1g662bhRW3HyQDAg9/DmJxUoIRjj3W9INLgz1tHJWRJJXkI0lJ6yDRKJlA4GqCztaf1rFFg
E0kqNZRC/QCDez5aNQe1aQvTTWO459fLnCO9FsQMOow3t2fA31MQmBnlWTLuJr/z1dZy7djq/neU
asx7UES0/Pqkyv0dQdTM/IgfDNl5/k1OSQS7fu8nxYbE9KvlAaZUPV9tqWKRrwhcfBg25nlkMVrC
q4VwDFeJB/rN/nWadQsoxfy3gDOIfaetbhfHoG8RR8yRofAE0kdINcYfBuJr3xfYmjeB9JxwhdNW
EyKwOs2ZbC7eGY2Et4eJ+BR+bWmXXUspU1ci8ciny3R+NpveABPE9aHW6eM1SRB5CcXOy1aGA3ug
rCQDlCgiUH55xYX+fkVNp8S0+bct5L5POMVvyq1rJouBbj8wSQLtMwHR9ppN+jtXivMoD+icX3h9
hCf5dAj4iiJSqQ+j4aXOB+41byFMhCuAhGjYCYbRHLiGHd7U/nbqOsRYCTpZWHiDZuPI62p0Zft6
3qlnyKNMB6280kdDfKd9oMRRwh58OXW4XF+EFO+5FJ0pHXrlFTZV++vbOX6rMENLXaK/38TkePj+
8BiOSpnTyMTlgW70LS4wwir88IVJoKvMSSFeWLz6TDJEx3KF1/xy9fLAIySJZE4v6b9LMdIBrKc6
QEj6cQnbm4FA73o2mn50FzhyeR26V6r8cXF+6RJFU14fZ7/eSJiJtKqFZJJ9mN2PC/CmGIziwLC6
SunXTaMShhipaTlrQgHYeI2UoVkbz8GC1Bs0d8fANUteh5i/85cYrs/Ep3VCnX1N7FMhhT2ahQC7
BGu9FKwX58V4a6N52KfEhmaYsB/TCrNmXmHHT6vwlyx8t4G0Mz8xK+SKPG8ODcF3aEY/0vhMQ7ZM
TSKwpI+/8ong4gpNgtTubk6pNOoxdcZ9T9iawXp7aY8reWuyfn6prG410D/AzOQbqmnXCrapYpO4
VIZVbIED7HBhNYewsV9NRGeWv5JDjRZU/C8OwWWFhUoYnndoxqsVLT6lnn9dN6KO/D0BDqkpBiYU
+MYBkQ31PSY7J7WwPYamQfU/kNv2ILQul8zWoEA47AQzR7WsrkPhlETPezqRDuHGZb5I8XJvx8Mb
9eSAx6cvxXBNHi6edT9NkzrCcrOTK/P/tGK9BhrAU0kP/CxjKdORilzMh/pm1Qn3e11tOm6MUpuK
pNbxjjQii01ZoBE9eKQSLOaqbOji/XnG/8yYU8R/40x7XJq5hYaFOwBN1FmgW+3ALlCj/ELCR1yW
P/JUtBQ3d6lJZ2i9n1plVxZRDffWr9vwe/lorEfMFEM7iMEeWSc1qqoNAOhMLOKqUWBg0F/ketJP
uveGCMa0gvcPz1u3MvFgB7kRQ3upAh1QQCFZtAjUJ9yLb/XzidCcMjzeMHVi9zvqbdK17EgP0S1n
m7vPWcRgCNOTSyzuaoCQc/9YGkkqGEZY2ceZCmmDMWbyP/B1inZD+mJW0Wm29KJPkuCbNp9Xmsly
i900ZI2d2oScs0gzxc87S+H9WHMCRde4VQTFEG3qq34hzTmM7S+Hrj2QwWuJ/MddF8rFcCO7MfKY
sWXqmO50MaFTsjRVKn32eS9u4D3bmFXFoebav/Hcu+//6ZwKFCxJTMeJC+Q5y31C+J0S14B1r/dZ
YegOeTX3ocLNoGdvumEHUvO6st3YXsZN51jQfEdEt/C3n5+ntgwgqBmTKPBV0qu8mamBhPkcC8mB
/oNI2hzLBkRLvZLl34Thv4rtpUrPcsRWL1R3DCldMUGkkJUMF6v9R8SKoWwPuMeas7uAKcIEq6lk
iGBK6YF7zMHx+BPQTDLOyVQtp+PRD3zP0lALZCQKKktjJQ6Q4r1XCsbKEXoFZHz1h7tV/M9d1kVY
NUluYwjVvNtklKjhVSMtNTvPVUlcm4BffTRA0US7H7lJOPo4Px6KojnpebUiizFTBGwH1rzy8nKU
Q47n3aTHagPM2qtwF8k2qe8TT1wOFB7cmCE9tm/eXVpiry/POJS4aOGXwaLwJuKn/pRpwqROU6ef
YtIRibRJqyOXJKTvEyWe6pa5YxHu8fCm5hqU2HxW569r6sSssAMHkoD98e6vJ6bGYTGQdUdzYBST
DkI9/+q56ZRMr5erEjo1DtuEyGCupQ9KLi4n44Olsmu8ukRCHI5r0qHiFcjZkfLjY2QmZOyMT04f
I5WVXSc8j4XB4N3EqZeguP9bqNxx9lSMI1K9dwb7nz+E5iifnCQzqAHPUgo2m9U9Im8u5DmekgRM
yeq/25avbgqgWdacYdYu1e2c00eEbtI1rVV7skAvmUnpkMf0r5KJH2C+tVQ0UHZZq5sMdwSvuzuM
kKFIjy3OnA6Iw2SXNrk9YPM067E3cJ1+WP9788bYaHbKsVmz651so8Ege6sGJit8aSwokK6o8jUL
T+TKLVp43azdt3Ht+LPnbQmlaXClZ+bOgrQywLSa0ONQSCYEgv6WCJ7TFlKA1NVT4br8rI0SkpjA
Dv2Xc4gpchkOC2xfrFV0t9t9Dj0dOdeMGDmG0z3fCUq0QotcUlaqHktQMLEuWbD6ExNZp0LYhBRh
WKo3DDz8XxzXoU5JFxjei9qztFkDdjWd6y5Sg7BjZHLlcnyKEyMkLqYUrmVw417X5clAB7pJlVdl
H1cAUnPb6vqUzq42FKI7GphTr/2G2IahqBTstlJs7q2N2DYXiQlHV3Q+T4JcyIV3OQ58QS4ACKXE
OcCHEiBwPd0zltyE7hBiHJC9Y190OxI5AbcW+/M086YXNkxLe8zFulH6hSlZNyK6F8bApTv3RiXe
PyyDeo4OIEvTiUsmg49rNAUKNwJrt84YfhfkKNA3LUQqL2lY0O4eCNAAS7wtR2Q3Shvuo7g7/Px2
9aMhh88xf7GM5MW0i99ezebFuwPb+nR8F+C6pHXpFnUTLP1z+Hd2jv7KA2CAIAmr65P9w3jcPJ4D
1h59UD/hHF/sU2WH+ZDrGnTRf80tjEuV3OrpxuZashElHP9lS8PbwGhIxkx/89YfdUA99nYPet2G
O72yq8GQPe33b2lEuxtHMiV/rAUVbs4Fmcl6wx5DjMLhDYSm7+yd9L3PIgGLl8sQJAUNrqDJ9MMv
0Cgg1I4IZA9kaGPA03Zo2LYk6LG2qKJBhDC51AsbTd7BoCNE0rbN2FeS+0+0aNLYhks4d5SUmm/0
uxgq0w26O7Dp1v0AnBlIJXKgfjP35UrrgkZv8aypqOY4wXho0EJmiFhIiNwgXbQfCSh5ffzFe4l5
lwP5l6jHv1oDbfoPSXcnQdav/mMVjOiIOAJA/b3htfeD9M3AD9UMimCqOHMCj3YCO19zVBcMbc4s
9I+OmRlCmsehmERX92V3kPyn9KVuvj/WS9mTJawEXAXbS3HHHVb3Ljyih5+gJHNHbnCh/LA6qMpJ
2rWjKJvCM5fPC0wYNTb6KTkfG+77KTxM3jiOFNRvAry2SOGp3PSbkC0aT4yA1+PnYcRM+0ZHxYZ7
wO2eRyL9vYaFgl8qx6elAMpp3nmG0zSOA1dLrAvuauKDsPKknInHy+bJcgBvEpK9mCJNWADNxIXJ
HVe9N/5vzrCpp7Eqxobwip1P+AWL+TEPHKssYRJd9zWRD/V5txaW5naetPXAlyr3ULlDdo0dTIBV
hHLwQBTIUao+NlFPpo/uiD6kH6e/TRXF/Ol2qLjTLz9sNVloY9JBvcbYRpEChAdpaW6/U9SEsHnN
eEqLB0tcJy+2IlASDnkA7TJUYqVHMTjp1reswCpQ1PI62C8U/4cXSnwo1ZpI33NsbTqIWX3g3Oa0
XXc6QHOJkYq6GOMJkBHVpgjno90Mr4NYCylcdn/WU8qHDXcEtMi581EAHPRkiQiibL2nvDQH1eOy
4EDDL1o7ZEs0OFHAy5Y7PRhddwio/LfGrcMth9bMF/qwFfbP95JrUamOJlrC+9I+nXST38BnpTGV
XrCJ3Nbamvroc3EyCuUR5KGj7jlt7a7kZBdC87+TB6qoHncOmLPVQCcbPaPBERq5wRyorVXod22P
WH0zbaWtFTn/wMS8hT2K8GFXYUeNef3XZebga8cf/S1olakoBf6TexPBhbHJMK766j6QrV6Yq8Qo
AqV3brJjPNv/+E1kT92TamECJm231ah4hNZ3KUkZIz2dAdgUgyPl7Y6ZN58CiBqS6ws8PDVMZJ5u
gjzSNp2uJmi3ZxGd2mEM8c5lxgUHkBYH9MXAhQ5fCW3cNb4fgmZjonT2MXlzVLpJlNmosIS8Ozka
pPsC8ytPNEwAWR7/SZqMkJaA82qyVPIe7KyjvxhvOdrx6ZUJEk/++duoNLgDIcIEDWSD7C8gW6C2
tuWL0mCmhi0yHyi9uT9Hcpibuz2DFdOm1LNdPg1v7WBu1AxmAz2/4L5F38Yj7PfaH3bHyU0mbEo1
1lZ0tlJLSo98W2JTMnoO/uxbJMXg6uB2Oq1cFeobZiKrlXbSdZOgEZTUJk43N0oLEHkLXQ4A0VvS
BukCkiN51g4w5TDOZhveaW/OBd9GSxv0EkfbSaQHAidyn9X3ki8MbsJ6bO/tvAehGDR7Dcz9PY+t
2Z0gPrLT1bkvW48bloZmbxJAnVtmJjzO2hmPRxVqJbUaa+NcHmwca6ZE4CSoTTLVwz4tooyh2HEC
yC69DV5PZsfDFRvEvh4miaY0qIvBX/wVVF8zUrgGI2NTA4qIeogvc57kTZLTVK/XBpR8i/P2jacK
2/T/HllCO2knJDPmpdiGwacnlMucJGDVwFY2s6QKF0S3q3/AQYu24tGVdQfH5/BcNSp670v2dWh7
HY//kSpAjpMtQQzi6HFpI3EL99gn7BXi6JSGJirwMoWzVhg06v42mEcDepHggNf8DO70git9cfAf
y0JduHJjTTxRPa07G/p1X23Va4cSs3EeD2YLEaXsLBzNY3/HWYMKZ88tteZr7+8KhFm7EMgMSLRa
zs6qtMuvVMovw5mGwwmJrXG6wC3ZoyfO/Q6jaVBh+4eXXvcMZbruuZCpgZdGI1J0M9OsOHYFOF9S
wZj9u+q+M0DhT0q0O3A4jpVRJ9aYkRSyvMyJDky12kKGYacnmveIBrYdkdqHaa7W5zKh3x7zeGGY
fwccS4WA7sexbhqzDNjbt7e6J6vmzLesY5tch9y8dYAoI2QQHTNSeDTz/nlCIhJ4Guycisv57x0E
wQW/r4bgX9jRFvcqwJuC5JoL5jFlXZL9FH1sb47zrImaaNsbhDedwWqQcaqbrWocp+dCZe3m6+Tg
paagZFgvrdlLomMl3Ganfwf6UCQY9BfPjDP47TiOO1MxZEJaOVDiEqE1g8wt4MiawipvhkHZDXoe
MUD1H14hkRS+HtOssrzc3G9HsXhxFYFW8KQCF/0AYHyegLJj+MvpbPX3JjgLc2j9aLbGgaTxkx6I
Mr6mczikRkx6uvtiEUJmzlWhfMY9nQb/R7xzJQ2iTiWa5kKm10WodeanXZlReDW+8SpqMFuToZQL
XQDnaLwEA/I6kED6KH9r/xLSuMwK+pVtu3t+OeoJ9ESdhbdBMsYKpcdyyAR1vZRCOCABdmLDrGds
SzMTw3YvLeFH1ciIxy8cbzgBpHKsQxHaBqVFn1NvJ0EyaFClz8hvOGIhC0hxhUQbTecIBT5xxepb
BrOA0nCtzRLXEoTCqU+AZVUc69bwvaBmDWua6r7ebRN746kpzrzUwpD6SaDYMP4MmI2OWRcX/9WX
NlY8t7y9b5NuK/72Ds4fIcpQsHupyet4AE1UJ1nalQW6GybBTOvEpqKwM9RNeJfU+tuSfPKU5HTy
xWqprvSgSxkOXNRzZWhoYc/sIhHjeSi4msOcy/8iGXL97tVZzmwLcmaeraTxkgyjae79YhEgj4V3
Wjyh5XIMj3J7gToekXbTbauJlUVCv6MDGC23MG/TZP5B1IdjlsOG208tSJbn0N+dTbD5fJHeTkph
7rLYMezmLc6J6rRQKs8hTKl7hoil3jJWTs2ZLbO2+LlC8Mc9C/pwCVSCrzDbsI7aDONK2/gnkrsG
jV79jL5JSJxo/gF2L2U6hW5FnwNvdRle2OOSNZdWQIP8nQF7YK4UN78xwTKVHbbkKiujCjCcB8p5
54/J7riSJRCd5b8W9h+0qNnbCwUz9dDulE0VI1PJc9yZMaPg1hiQem5c3l4PZ3OsiRg4ynvjqMFU
5RwXwVU3ytWuTi3uWRrk0stW2cu8ZBAKjS5GEgopmZFhu7DhKuKFHduexfwPmf6KyQ6ngqumMXM4
+wdTtMyMUjQGNEBdrH5b3sAvlO7dn++Ayamvo6IIKtt8sUJDumZWaDR+LOnxCLetQWuCCybC0s3b
6jt6vEYa+XEoUF1daWYr+e4CRv07xACBsUpTkVz1//CTaA5ZmJs+cyjLBwjnPmN3Q4nb3iVS6EPB
hvPcRE5eW754jwF7uPrOAsp1al2SHgTfRtbW3Af4RHAo7DGp7qXwMKv/j3RTra1NecL1Ao0bYbNf
cd8x6ZNlzb/P7gIDYeEoNlFEZqD7URggeXrOKaznxVnpuIBzdn2amnG6zJh/cqeMFZfI/lm7llG0
ou0/oVv/LW+NplYeOJfSnqpgnHKM+1ciXc9f3iYC2+RpfW+tlFjZOdz0DrzXIXH072S6hgmAdr3T
KJ8wl/T/vrjHvnR6jIWiGNTqWbHaoH5FN75ht5f3QxXPVWcwZgj17XPH1MAl8IP4isKoRaAtaT7T
V5usimz/tl5k1vmPhITct2Ip/H0hqhKTcvch7IBBnDUCrNvMOO62vHLDyQAnK98pzaKc3dwf15i8
JBi2hWvJKfgAsGF9oA+oVPgplExJ5gd7f1YLBe0jkNpGdGwwuuq2LtrsNVFPUb3GkPtV9ypeArDM
NNkW64YKW7et/484zfFG548+JK4UPfe/a59FQLJ29JPrOnfg+Xar6MEz4g1puWjYBWiCAHwpvKsM
gn62SRZHR49dWmYRFKgz7Hpky9ce1rO7QztV1vMzSQDNS2Z2H2k6wa4+IRQ6X46mKdd9hRm0sbyu
L3GH7cBn+Gy1b+IPj5xdHbkEooN9P+SrthSASnMOW+ucqURSc6jYd4uKfY+IgHLyRa20Ap9EfVb5
zP3p4VVV18ZqIf4P8Qi+YKu3MIn5FAoH9rmCd6cvTYq1ACVIKTNNRkGpaOk09FeU3KYQ32nDfS7T
gR/mBYfTDsgMPxEO73Lew7CVrmM1NRLJZhGndaXin4+O3OWpf5m9yiiOtSraFb5feAhgBMETODqr
2qw6DbE94ojwF51mrASKRYP/MsyTpCSnArP3UhEgnHAEQcTfrbk7H5GrCGJltVcXH48IhUce9rCi
JHZ8jEWj1OlQb3tL7rLmW8mon4+zkNnqB2NGCARFsJORgFK2ks6OZCJnQzt09UhMosMZUENVd7Z/
4lfVXw1QCh7n82shr0+QMtFP1ABY5l8HKwGMfcoxKgsM5yi2kJBPu1Rb553TB+JurmaYpqRuBiK5
fzitvMfIAeosgcbLtj0hYMWsNSKXeWWht6Ax/9zbddL8BTldId2nRurhEP1pwNddiSFJeYJZjRZw
K6hX3eNGzg+XxNaDh9ZOE75Wnd/tax3msn/w1DVck0ZgKHItu9a7hQMCfQQvIZN4cNBVAOSUMAXt
l9pJ2QwYVc1MA53MeXgEfAsv/pKX0lKtxjZt/Gc91o71mAlXGg0/UfsGQLT0Y41+2E00ExS4wby5
8/fbunbO7g5cstKNl5yYKSmVUwQ1WaTTcClk1eUCU7icHEtPOazI+EiakCqh6E2OOrp/JKMaUtJ6
o0Ju6fW4WKZQMJ0D4ljWxnQLrCxZIZN8ODRAvN7r3WVFH16Xj2mty0gHCmhNci8xa01WmYSqwMGD
QhzvnXSiRQoFnYESGJaSjoaZwmL+FkvWu03kCt7WyvvSxE1yUFCOVptbunHMA9csNetRsLquLPBt
qhZDdzYuEaF/Aa9kC7hDDPaRqg8PpuZ1/B6/EaH4kI2GEy9wsM5Chw85lS34z4v4UDjR08se60FZ
DNO/mSdgPsn+wxUb47smY3VLZ9UdMiQ9B+iQMUCYkfz92sXD7IOBCplYia8x6Ea+V9wlHaSTIt8g
9NSeN5P+oYD7IMCaQVrSxlEjilLXsRxuUGFD3nr0u99swQjZkF2t9gRcjRm3EntFsBK7eM2ytyou
lFobXEADiwYsV6zPgW+wtyATl0qsWNSLWSZhuxrVm2+uweEfLXyqNsUHTGvPL++fE+WW8+iSG8vx
Fv3IyCJUu1XfPM77NKmrlPGPtGeQDSl6YJxDGR2tCbzFcw5p9NM2A6tOXICm53PeytLAPIhlNuqW
6Mx+3wILD8j1yzZvcjmCieDoCAHtMF/CbgN59GMS0vWF+IbWpcu9GlhxjQ/TEhlJHX98OR1g0tJq
fp2ZbF134Ab5mEpoNsOw1IpwoL7j09/gcBJdtt6490H3LoiGUWxFC/U1XN3yHpj+QJM+qIPi9n0N
x+5IHKk16y0Cw+/ruwLqcHNVH9MrJ59EoEo5qzA32byQYBfkTW8Yu+U6fwk7T5AlDXpAYln7jedt
uGAbmGH1PxGnFKUVCBjXYjVCwXvoCzwwoe1c5l849AI/J3DfSGb7/3KAFP+pfxzUHKwdyjpfjOTk
6c6QlDMxjKFwQiv3lqm7w5DrZ71cxlQdWwnYWHvy3Rh0Z991gz+joKzYIptXHnYGqLbC5vLAnCqZ
wB3YIjZY+4qaWYJPjNorqswxVo54V/0sQeHozSgmHhvTCYVXWW5HERzR4XEcfPp5EvPMBFC3r1eT
i+kvVF9sFhkzaOlObbKhyG3+u7g6yAE4x1PXyXbKbIcg18Xc6+FiR4TWPyvEfF54DkQ5xu6Qa9kR
bkdmmWJKXpvd1quqjTvurkhINBzQLIuDtQEk9Ui7EQJ91+KLV5pqhkQH8+6ajBaBXaosocbHCsIh
fKq6J0sn3SvgCiInOEI3g1uzy5kpkXeZJ4R4G0QCX6EdiwuataHkDHk0p4imVl/AQBx1tcK2mc+n
iUNKUFulDVdOVRUrTFYlh83ZlQICvo1lTaarhiNOYNHQ/NQTYS2NoT0vqXBFIdqWmyH1wRNqa6hn
NCgCW6klhvKo+JbKpmN21MuhWN29prKonBhzGASx+KXQFtNKSrLbWKQxUg6mIQzFw6LQOlLv1pAY
KhlK/O9doHU2lBObTyysWabG4Y4gvqWLFAWuQc+u96z9wxqSxqDmWnm0CHiFLAgjkdJL7AaQEQ4m
EDwdKYjn9Owwr7U9HBAV6+inXu2pecrBj5H/o4JepJSKwHAjYQnCF9gjAAgzD30xYRKFflaFG9tR
oVfqI8xaJezvO2dUfb2QYYFHNL5eF8TF0mPUI8n/jTqN3JFWn5/2vo07vGkeg+lMGAVLnbn4lcNe
cba3eyoV1y5wl9mc/fxOK6pJCDWGqtvY5kJ3YYZxgh2tga6WnasUBnQnx6mz+kCOayCF7/p3w7n+
nFPF7ThHPeOWLk8tjGnVZ02VpwA42y5INxuv75z50vExBWvdXOZ8M1saME5oWcMJUS5ESTqAN34a
BaHneng4oRu4N6eNpL7alT3x6gz6P0tphD3einz1IAfgQJl2DF9O33HbHmurQygl5y++hwqQ9XKB
oCYTAB6fgT+dYEhCpsAnFBTPHCEw7M9TC32PoY3NBR5efPpFFHCw46zQLBiRaDGemi7WHXAdT8Xs
kO7IWiBj9Mz3RQGAlocrEvyed0Z0Q18YbfajFXjV9KTh6QZM/aUHENpCZPu8fwrguNHjcEYQRNue
tvtuawyEYk5B6Knt7bwxY10ijeFzpA8mKuCOKz97rntLXMHGM/6YQawY2ujY+rrPAjO8kG407AI2
ieaarnXgvsYdT4s7qy9CX4D/2zLHTGGjdCwsrv0IoRh+MzoJvR1pebTF+EQS2fuvkdAzmScCtgKP
vLr2KcvAEXUyp0TbPc/LIWsojiWsRpcwiINEb+BuBVErmMB866DRLEPXGvfWNaFjV6ohNoWCza/a
3U/5Mf+ApYEQBMJif2RzXi4YyAeaWatImlVQW9Dj8ukDbKWo/tWvpGpHs0BeVQ8708b/bDdCFBhz
3bpqXxz2R+HefbHRCBkM/Tofs3+eJwjEoc51FQJ/epfG2MvQMfu+DCktNjItIalw2vMtB5I2tIQO
DlcLKp6IKgS74bxE4eUslY4Ckl5iXtwfkbIhJPexScEYeUTXzM2RV0xC9wpvJEGV34siO9aO/7MR
16I+DBuUY+ffpOZxsL9gmaW6bVevK/w9CcUb5VwnaEkCAJbdgCPT4HP+3+daUDLv+blHNli3ff3d
Xne6WIN07Ck41V28q3HXxrDguAWimRThlOjk+AYf+rcO4N4KrkK+YZSOKuP4hC/zYGzi1R3DAVMp
k6ga1hwX2Bdi3I6IYriLQ8m/EHqWe8TdRfWjt4yngvpi5P1JQNnOLS1yzHGcKZD90UnLk0ie4MqF
ydFFqyTlWA8Na0b+OAlTNJEFVgDI+jcc8an3syn49aD6tIA5dzodE72YYAKLMgXMuTj9H4WzUgq4
s6Fgyhhn1wOCxwwQwwFdmBcq7vlUOFd2KeaSuceruZFh69WmmG0QBK6tHnVQXZlpbEKFuChy8fvr
8Ms+IBOueiToW12k3qcPcOl3Q9bQ1kb8yFkzbI/5kRTopYMxFo+6QlETHhxgz5w3Nh2BR8G5+q2k
jenjMXA72ZzAx5OBBcN4vpHKVF/rTOwxHnvzkqlzd3dQlhHtm9WcksU09XvrFLaM4g8xubTHFqOP
p8a7m7qkNOBmkZl8Th8XwydE243x5zNqsaWOsV2LLfETGilreK9VDg2i2btJE47lRt1qBPr6hdif
S8VHqLVf/59d+x0o6MGOjP0yalO24JBFrpCO8zWa8ilHX58whbmXFT383PjzURoRICtMkSQQThQV
pemwlsi6jO0eMwos5Dp342bpGaVVJMrTDPR3e+bsPC0ssuWds8sjC8QmVC2Ffu23CvJ9A5WwwcYq
gvfNIbYzgjaIbODRlEDC9hgnaiqAuaOON6wVg+XMH0ybU6OHgC0VyLbTQ4saw7GBWE3K20LvPXCh
sv4tXSZiWYvxttngGHrCU4Mk7rMEq7ZqdvUpbeMdYSiBMKFjP+T2Wg175xx4ttVwPdv7cdXeeUPt
Xv24UOX8mA1GgF6nUpyf/H0GpgQtljWzut7QnPd7V6MMp+M1L92h6X+804gYequCETs+CBWY1g+L
fI4rBrGQHuzppLZPK/oN3yV5FAnbCC9MPbCN3dyUuKRNzioAIRoUxrZgOKEFYMNvT7sgQr6Xtg8Z
zsY9ghjA7uf59rVfT/F+LEuHB3D6JsyhndNFc9RywQE2KA7qbMlO7KhIyLr2itp04yqKPioYeJqa
UsoYvZHzKdmsfpsT6wouo1N9cpTLS2mozaZNSLd9PyqLemj2tyeVH88fqPegqRZZGnMsXRKsPS0o
w8YDlT2o/eekwcVzk0ez4JBHKh4AOYVliU0faa+gXQQzd8AMtj5yoOKvYMVxNtZBEB7qkvOt8RcN
A1gHzfufwsb2ka1xqrWWh0e9ogK6p3WGXiU0b3yjO57inCmN/WFKN+sqe4fxTHF6elkEhurZd2zc
dykLXTF9+1KoWS19cM915apC4Bd6WPlAHw6ECB4oZak4zBYeBnJKjUOhvdxCYK6cFnMOWl+CLRO/
gBBmGonyE2mULk2uucDg0dM5xyEj7NFl4JZFPWJFm0Tuh5tAYi93dbasmNoxyiAtf450w/SoLNop
bLr1seEibEmvftHg5enAH6/IlN7n4afhz/1MIumYcrQhXc1FxHZxwDSa9hHB7S6K8L98tXeM47+A
bxDWLpd1y1G2uvDxhYBaLSx83vWSDnFnEfwKqhiXXkB+MccGH9ZlSNKrZQ5aiwzSyWUQX6UMUWtA
6lkHIJh0gO2uH2otZMMBGxIgU40VpBXEu1dWOnA7/zZUEUXOOICWXs3xy9bwstYyDNg7nhAiuHBh
oK3gojBR+J+1pcXG0/I2cUuJXggUOM1DUuv1p9GOBg6qxlEDJBBbdPjQ4i1j0kyDHY3kT0jnug7V
imYhJygtu3iBo52Wr1gBDlZadiVxNaJan7SkuHny+g6H3gb+nYA90W3jm9TLG9d3y9MkngUJOAoY
73YCj5liBnr+/lBQpD4i7N5HHOsdae0iPQtAmETCq4kmDmNl8bbCjpYHu+gYxaMKO2yLhZNRJiaB
LxdvtVBpW6uYPVAGHNqHgvZ8tCK4xHFa0tEJBdsLZKQWeg6QxxqTXU+Rl/lTTdp7n9ZSNiXjaj7w
uq6hZqqFWvC0qJNcjiKL/j5bLCASk7W00IzokdHt4KUJFaPlWz4gb9mnGGNt+jDmL3/JFmdSoyoS
HeypDZ7UZk3EX9Iobln2lQAte4eS8o+idZ5I0baN77E7lgsS8GumFlFBz/YZZKk7OkqtC9bmYRc3
NI5m7vP/m71LDDCfZglEaH2TEA3wPU0kONAXBQ3SXvUkfV5Fl7+Bo4w7CyFvSDxhdvMdiU7hObMw
4ilirqyzPRtCW0eQWDj1DmvUpk4VEtTa6L32EqwhtTLWYZL2YX+DZnsw+ECy5nI9FdSTIhEsw8hN
rVbO9PRGQxeLbwfbxu/oesf75VsnJKzpjI/mxNh4zJ3yEu1H4UnhgtB3ODRdvhY/I9PrGCx6+HcC
6SNzR6xwhrLXfhZUi/X9H0TNwPUdVqTxeJDCf4iNztFlifQmS98wr21JOMwQNqgIXhzQI6LewXdT
50oo2BhiHe/6i/2YvAKT/ufj98W4lMy+rfNwybu/yU2g6rblQaAfOgdIThI5kQQY1BYchGJCfsg3
BQXAHi9R5xhxNbcTko+uouw3c6bvFuseFP5tbfg3AjFv8pnE3zLEHhDzQkBvt+5LsfKezWDeHKkP
dOlYfPYrULwNFT/iXMKYKkey09rzLO5E+QqAIpAm04bD8U15cR0AtI9YDwkPeuaB7OxM80VtNp4W
7nk+nwn85v4ek4WwvxXSR7WXen4/J2h0Xi5cbHn7fmzup8gjKjP0XezK+vCxFcLW9m9zR19tdKIA
ar8mlErQoeuqcRI1evhTAU27M+HkcdCvypJu0SGPmwyyxOdgQTEcIMi1NsGni8IKZvQCH3mbWHjG
PipAzpUxR72RSxP/9fyNS37kaqRnnsQMt63FEFT0RqwwMuW3h6O9OkHRpkOrqNqKNC8dwMeWoMHe
u/Q4nXdTYFKZR1947herpozSfi08k9aphvyadjUr9bAY/De3iuQGI3NJrWJW5TmsVoQLWQxtQipg
TrLqn+OEa82j67ma9T3eMi7QSoOY8nBs9WPbrMX9LwJB1kBvQ4kEZRauEXX5RJJuYk2dQkhx8UZB
fezGZus2gZWZSZi6RIZyzi9dmF6zQmqIImAxS66qtV5EUy6IdjPJ6HjYmBf7+VIqCYkLdEQL8Lpv
kR9ytkDnl6wjxZiBKkbMN6k0CmXViYkKXYSgWdNh0dgLW48MK8Ly7p3++TfCp2AXz8TX83EgpewA
mnlG3jyIPlIdM6RnYTZfUzyeqD978xgscCbYfujXv7vVxoktXPtLHU3a93RgVyPowHIEtrJvnXjw
uukf+lDoyTLyRZfsVAHTlUvDJyYN7hgrMM79aY8IdZhUnaDBbuag7CGHovqEPZxb6zfOnhOQCG25
oKTXDCYxeElBHgi6S/txW7fobefWn1F5IzcUvin6V9ZvjijBlj+joR0NlnBGsHVZ8ae4xlNPlyAZ
tbojVdtaVINanLA98o/c6kW4I0N1kt81SZKqcngCdMw1Qi/aYsfXLMMMzeij77CSgi8hsTSMdWB2
GqnO/le08ByfuHg1uac3RS+/EwzbrF+KaODVSRBNHztrwDKL1nEbGg+pMl2kzvWhi8guxWT1xsrw
zIMt8mfeweYDoS4XiKARMt3Rn2XxTZozmGswi30uP6JrFZe07XVvrC1j4j8tFBsRTyQF+vOwLjw3
XTfR0DsA5oKLYlqhc9hBGfWF1r2jj2NRp992rOrAcNpXlZCbPcGQ+d9g0bd5RVQnuBGEtqUDwf1f
q7GOFv1DyDtG81OcQKnLaVHURgvZEG4bMj7J36RXdHyoDE0BdJaC8GU7sj4mj/ElM1FVKlm0EUm2
8q0Snxxi2q0Oxz1hAcWVLJUFLwEk5AwFvkGOWmfhGuebqQ2/MguXlsppKnStNG8g9vRGt+2Z/r+z
PymXdaTDXhh+rXD8TNPP9Ttfxay5vbDcxNVavb4O6N5a3Tz6RuL/97mhulpQ6UYHH+4Hqgx6n34o
O6tPX8rMBXHceLbp3ZkDCsv+srfYQO47XHocCaaALicqYSwBLqt1N7ySY3eObZy1V0XQT1wn8tlv
CgYSERK+ZO4oYxAzCA1MAnGqPCZ9W4Ezvf1m+XoOMyvXVO5HjuDbCNvBFGqM+wgsjLPBaGytMnEN
HiXPuFCQiIfMUNPPQg/O+mI4shLxkcDoiJjuLKCQc5buq4KWfHIO8TvDGRV1Le06PJe9gYWqxjk7
Me6vYDQACHWFzQRoOwyLbv+fMQKQIx/Pwp5puGtsewCjaBGcwBPmfB2gOxydFvCHmCJG1/6IUSj3
fmrbz5Mu/bsgiVSaE7gVMc8NOgFjXJe/BTQhJdQZUW7dVmXpxtmKqK3ZN6RBRnadP4IPINaTOo3H
hxRmxkizNj70ImdLIc1YBrNerKP6O+vPWAZyBhaFqtdW7EhJti4WvLQ2PAoGj0zXnaHdMmq2TNXX
/er3/3gCsYK3vl1FbLJkSzs569c4XfOvvW1cCoM3NXHLL9ndrLxPb43h7kpft3Z1/ycfm6P1Di6x
QkVtb8CJdQaTWq1CIr/9p7iGK53mEAr+UO8PSzU9Mqsfj5ZGSDuNZ3686RiOm/vOntlB+ZTkZRkE
AMLmbc5ZDWCr2062wQGuYmRfyXcT6F+1jjI4DoYtGW7xMfPLbpWjKv8Xv2Q9kYdv7YceKl6SHiNT
98t0+N+TsCg42VSchzHIQssvh5GpEFHNsyTujzCWLIx35kXRtN5YmddssLv0yWZDQ5HH9oLHB0Ot
5otbXgoCoyiWvy+4MedcqnNfc63IqXvcfF8oPZJbspz9o65p95g4tlHh8dyy6jrecSH0xxNXPb1/
ZPUEPPwaDSDd5zFalcgaG45Xnn7g1RhxQnFvM454UlOKq9q1Z/vd0Cu9ouFhAUWl9Be/P0LZpUDD
zIOjq3fidDUPRX74Ra3keeMzna8wXiOlvon+H2x/W+1bFQ4GnYrc/JFrkRg/q+cwdye2NOrb5u1j
GxvadgNAcREbUWBMYSe2g1lksp/aKy9146IKDik5B0LsILmBc7l46P7FCow9jAlUqLNWP4uCVgN/
GDXu+CF1MGgAAeoAZvLlLNuIHvS+dijcH2rEPUp3XS8siIPPcW5N/wWmxedA0DFTLT+yIMn5b2/7
lixlDetNH+SSyauoWhilT+bOJQaj2UadpCAqWvij0QN4zmKn1O4NOQjGjKj+5su6verxbl/YoPVe
lFNC4TdxWx5ZuIUFW3rpUvUjNVfGlqAq5g1H+jHFhfQdd9J8n3e6pkp0PD8R0AHn7562+WcTrj6f
9bgdftisk4bfaGkOKP/IqFSXkb8e9hGe6HJiscvAxIwA76cjb27/UN/0Nx66Fy0wSmIcN581o6Eg
0kAWdanVSBodiRhGCdF0O5raDe19lI/NKmE9rHFIWOucxkvfwvVkXGATpQa3A+JjOewIEtS2q+ii
GbN+/O0qpmJciMmiftZeKG0NrN40vlBOH50KVopGtUgpW5N3xAJyiBdfUyK/hmsKA+0oDXKSx60H
Dd0stWEW3AUbSsDP4qSY/Fn7I2YNbn7yhybis+ZqT7NlevRM7pCeKPclJCVFm2chduR/3FvQPa+l
lx8IJ5xe61NS1+SzF3OHd02mJrskD+Dp66gVYSHtiDSwpAeyKwfEmx32zpHLqltLt81lIoAiTJZW
WffW1VjdCuihHTQ7Pwyw+n9i/5+8WUrCaXPyKhou2fTl4B98/kKRzzS+GX5MzGF22ZK4q/Pa0wPp
73omwO4sMy0++qMfikK+cpU69y3NrJoeefFWJfD+4uiTTydAcJJo5tGxAfEjG4Jo+Els08MdOn6C
yREQzIsAOLARi3MJ+EOfcg7es9rda2ATVLZ1mhlKmR9jERLLG+Y3IR1QyhFFoML0a7ESr7LJ3Tck
tiNy0iEmkBRhG8y1YN1NDmsNfa6YwbRKxBiK/pU3tP15yzKAnFnSxlrjGJpEWC1XXbgVvfGkGACj
jI1dYX+clHe4PIYWyDGCHtl1ow5iqYDIqP+eIb1E4zs9x3lFqDBMVir4deuLLzVi5E5n7JHPLGHq
ILATyUNqjRraxv9jVKT05730TrXjfE3ZeX2j1yMuy4jVkKbaQjPGGYDDt6yZ1wD7IEOCFPm+eqtY
Iw42M6UhTtNvHWwFdksq4opQqXKhp70ucSm7SbTMhOpA53BQ2BuqssbV/X9k+HLg34GEA746Qdni
ayH5RYFn+gipyVZZ5sGcUKDXxRAF/VAURDdioj8lLJYwjEYsws6IGIADdl383s+2SsdQmwbmgn2F
YCdPXKyLrnGGPKYxdYAgo5KV+3GlGOneNUo+mbp9phJnTlK5aG5/ROhCeGDy114O4G1NMTuS+5PH
KIwsUcRlgT8VIUoklSUP1MdaMMDDwp9u7chWtZDgAR7WF+Qs1MbZEJQyfg1YVsIK0FjcPeMApsAa
8FLQhUzpAgjLEXN35oN0zoHtr7MEGsRKRl2BNpkxwRqDev28y+8hrdApnET+sgfNlCc0TGfFHtJT
4mspavAWVefHjO4oBhpCQWPKcUPhcsAAXfg8DvJ3Id1FHQXc1jFUq96gkbQK3LBojUNgFg4ZvaA6
jLOVrAcYQbu2idT33r3o9GSFculderXgdvOkXVESf5dPceB3piForg6c0bRpT0oC2OFo+oTvlEdq
xExSwt1fGdcD6iAyZ9fYqm1puKtwU7MfL0IM+WrZBLkcgg9Cb8QYCVd7EFCICZnVcYcJNF4yMcA6
o/b52wJlNCWyV09qC1TA+xGXUahaTCfE3NBQ1SzZ5lmMvyKPsotzOFR1BgAupGsw0LbW52Jsdajp
L5L8xZ865QjF8jel1kt6QdAiHZyloEOjG5ewoZRvJuYlt56H4ysPXlUq9XDHv9GTbY4zVsONaig3
ksWtggZvCGd4n6dr80OzEz4bD2ih0nIjU6n98nWtpMAFyqD+23/e/UYQl+5wqpO+LT8ouBOOuT7K
al+hQTXItQhJQvr1UlqgxDW6VKOoB0cnD9tCXWBMug7N8VOBg+jsdl5K1iyJ76wM+IATpC+9QW/U
evUUi/rFM/axiw6dGyfnXeUVoiBK4/chR51lSgJb7sVJZGrNk/xPj9vDz2YEtPp8yokZI9ch08Yf
E0P16uK/TBWQVfr9A1c4V+d36/+14y6bkkvQe1FsJWzZjKZAFkAJ51nf79HrDCeMhVS4sgLqT5ON
DcmXc8xoDj4uiPKHJGVOPoiOLZpr+TruLrJkyI6gDRr9n1TH+xRy1DXrirCJ9Cvv/oStYJsfQDE5
S2CWpHNm1YXqgXvmxvTFx3OwWu8Tbhd/4Ndaq6x9I2mbPQZo6CMinv1LbGbW3beKLHPW+cMF8fJp
KIiqccOkclWAfQoDcoBk8VZEz10cJ+Hfnr65QnXsHLgXG/ecQa5LKbnQPSEYQMp6MYV9X0x211cG
y11dB6fTpSO3kAYLLy0iU4p1694GM8Xqdg4hYE+GdCtnnQZxru1KjucXHWN1SD6fTDYrJV978AwR
DRcLHEVS8p4BbKbiJwnpeollu1lX6vWdVU4wR1VuGwl9nkA7iw9/FSAAsCx23yM9GJHYqLLI5Hz6
7acmIOCmxRjEA67F1f2VqKjGdZf2wuprlPLMA3Oze5zt6Tf6CZ9icxETlgmYZPeRqM0P7gRgeYsl
M31u9c5xTuGwHBQUJivQH19how1uHOoDWDZRmbram24jUBYZGQNaLrtybVx4UDmC21eF2sWqGfPN
0MZHbytWa7vXpdsZZAx8M61GJQUxFvrFAo/QZhqs3qV1iqJTem3UEegvXon9QeTEdX6781nWvfdw
s8mEge3p/HHfvAejK0t2zOy7Oni5qmv2IqhVXk4vFmLeDgcTj5He+glZGje9zCR898j9axi9spL7
kMOo96TuNplanmRLfode4teS4FVRWSxEih3xMV3GEZ62hYcbdrbBj52FGwjRDGIUM56wBs4fNL9Y
8gWkIOdPst0AlkAhsRDjedhuqaXqbqYZrH9ACz185JmUh/sGD7TGkWRmBOFGGefv04oPtbs7Zt9S
qZYl4H4sdjizHEpnHv7kYVJNDxVsmm6jg/qTbWLtJ3CwtA9VN8aTUk+7sOwUGfhSGBOfQX0RgPfg
dgvfD27tsWYsLYdTLEEVGMXoS4Em+6I5ymlDgxf6q80SpOOwF1sT5k5toSpNq7yolMdQ1tw5ZN2Z
sorcgpYjK9SDxZFgciFBKPKB4diEdwsLFmk0LBb16Xu3tsJ9xrLylz68Zo8sKA/Q4x2gEZIJD384
GrBRI5ScSvEs1dUcCtiLCd2IPSgoryseR+5q958jdLpesHaDABjhitLD3QpUKz/bp6ry98Nqk7vA
QV646ClJGWAOsD88DZg2yb0E0W9ZVjPTzXJaYgxbqKR4707XMYBGlptKK29K3Q7FWlimQh4qIDiB
ILsV4JrEih+9zQkUvd7R2+V5E0GJodmlcGIqlLwU/x2R+Z4NrWHljRXSi+MQ+YKpizgtf+Kwlw+5
vxBxpzEYb0iRqedgSVFfVG6g/XhA77bW0yUkBVv/iy5HfjFhDoYh2Tfk+4cVwa9O67D65lBvnGjM
6kjHqMHu3FeGoyoitnPAebxtnOC4m6k4P/pdscmLLrZx//Wqyg/RG/SMDVo78zh8CUgmQCfXBKoO
fVwVbEHOqz/WH8AJJDKh5Df6OtqNgeoZ+ZJMTLTRizrsnhDi2CdinbY45ETCpV7QNVc+0yV6Unzt
kuoNlF66rFsahQJYfX73k9GSGQucETY8Il7UvNAzWo90yKTJe4/x9n2r03cjPEOVG0TBQEL7G8h3
WNgtjv91dSjzAEnOzMaZHBI2ZyoQI2w8jvHBq087cckt8GWXVMFGhJGGPIUZSVbiMdEppLhrnd27
as3Si9Ex4xnQRj248CYRRn/LDomwuKaA3fzI5OrDmT3SSDHN6X8J/NhZnBAxTvLdVgJ/anebwejd
fef1uymCVOm572EpC2XGklnUDzHYcsIGojw+UNCjA+spEjh75s2XF8G6HjQZuyesTcBy+M8ka9YL
H05As8vTAqTBylESDdn4gJUibK+L9rinoeMYnOY+3s9f3LgcVfRVCC9O7gBlUdWM6nk/kwIsV1Jq
G8UunMizVIoMT7Umamh7RMOKrL2TFDsKzk5Y7j36Ca1Wrc0AwUKNaZwAyQ1pPWOthE71RFZBDs4S
UXSzrVJyrebTvVQqdE2AYccIa9CHyE1WEo/o9XzREvEqn2G68JhMsR9s5HymIL7/YtFaQfcOoWuV
LjFS/Qigt3BxJJrkPP/UptqDEdzAE0aZ4Zt7aSFaMlDb3uZSYjRshywM4TTJdyMwozToL+Al6//D
yDXxdmwfGsRnNHzBjE2KGsvo7dXHwmHKHVWre0pfjarxzrW9QhUPv8nfpb76hfyFLpMVKNrP4ZCz
WjrgVwqs4UmOfMwdaDyexrWTJmaG04qL8Mp8GcosSWEwJ/Rjq1wU5MTQB1LLIAfEljjG2a6TLsQn
7mXzvgqra7tDp98F/ynsIEqVvcWQV80BJfIDDpFsj6Lv+apBc6jjnjeKhWO56z2Jf0dAp4i81H1r
4AWdvvzsc95Ci0byvIToWN3XWRJlAURhA10KJmB34N1GRuEAwOPCLJJLmRa6Un2+Z5q1qsK1zo4V
SFIbPBe5xoSHluHcn/M44xEKwMFT1v3rnpjQXYyebO5BG2kEKvDCJKMLSqsPa2JDThzrpvwVeFl2
p4gVpv04KyGRiUnyiFl4iBG1erNKdFSAV9+5D6AmuYMrCl360FSJAKfsLQ6BC2ttjA9Pvts56USj
HjuUL9uNWDRVj8+K9CiAp7aNhKiU+GBiXdFHCtJ6pIvaoqq4nZMaBeqpSui+4aVcZ/LSqx1ZyF5/
uiDkYt4LLFh7tMFMlKNGg3vTHlZEDNDSCTJDdYmfjpmpuKI42lHF89zWnZT8Z1tcDZGxfGg0ZBe2
qRCgPIY2kDp1md8yIoL3xrvnUGjkL9sntRYtjEDgrFnUwiL+EzAyY3UN9Ioy6TgZjOGFrZgRZu7i
4PNYxjJpxMJPlAf/Iip4HDNEnogqiv5uGodiUwXlnLcG+3NRfcXh2MekWoNT/KNawzbOd3RFnO82
YoEpdgS4sZjTVvIb7JhQTJRtnz8tOUp5NZOYnbDF2Oiq1Ck0zawO1G3neX7dhLO7yJZkuk6f/OAn
O53mPa9UpxQ9KD0Zk/4nHVfY4O4QvWQbK1QWUOJhLQ2Csycx5qDNxk4jnbT3Twl0dsqnRYEVZJpF
7XzEPYUj3RfQfclg+SSp9PhFIPaYG0/rjn5DkbPCxyDfBtHwm7ibSEBKq3Tf/DLxV8s1R1e8D6Zv
WeWxTHfgIvm3YIp2MKKzKqKNhMpUWvWZHCRGXr+MV0zp8pyjLIc+ab3SC92Ojei/x+kF2eMXcBvw
0F7zIQDgbWhlgDcMIOdaqO4Q0XhqppaHxDCobOG3O+MYkpqVqTWHdEqoEwNZ3ZRtgMHnxpgzLJSJ
sazrQ9cppZVS2+8mAsZKZg33LPz3ynB5oCYa4lpnO7Eum09O+pHLTuq9mqVXWW+w9TIDTC4uQ59t
cRHGXUH48q5/8hjA1iTvS2jTR8Qz496kw0bfVlTlnxsTzNDpOCAamPYQxecrZUux1ED77sQzAYQz
yYvM4TFBjBD4R8S5AbCCIJhrxrCIErjhKCh+9mIYLvmYR+pQCE02OQhPPLsqYpODXiDhUVuTMpIj
qm4CduaDhdZfFjAKbqkbgFrE38JL3MPFHYNLLNTcALmpTgTZgLIMomCgBFH9YXPK0JhtuZuubFr6
8irSc52A/vC8tco2dSBLpjoeux+j7FeorHCnaJTSkxfMaP8NZW4qW/byHH63a+iTIUOSbrMA8slo
FaTChBXiZsiekTTkV0qOgukGSiqMgh68LjcJWybmQMYtaYDxsbmk48Qs8CehSu1o4Sv1sXo4W3Xv
b7LNAGoWRc/OAfQqhIHci4ztrezSC46RHTqe8YKIfCK89sqj81fBBOHYaKVhlttqVsBonNaFUako
EBMaYFW29YqIEOSz4P4ocqDykElPoD+ekg8cMI8pHbonx5a6xGAgrfeBIQZeztm81J73ik1NWSDg
trJfHPVuXQJ+MdJpTUZMA2NM3Eu5MeZKz2xTKmran8zfzfzpZbKkQMwMIWS5cmF7MRJuWWnR49W9
URAKFIUT3JtwyHTfeiOKf/GoRPKFBKFaSwaBFLIig/ueNyu3Kg6TJZXXmmNoIVqfnnQMY90SK8zX
LhvxRcmPBwYjXvf3/dBFkyiBC26rTI5gGfeADypr5Bc/AzttMQcYCDRKkkp84KI4eoPkT1U0vby/
ybxulIlCCp/68TOG5h6hDoNvWL5YeceIh2xZjAVMLa8wJUsQAfMJC1V+hkiZMECDaxSbK/rnBOu7
6okDj/HRXhRk3x/XJPxKbmJniRWU6+JsFIwKu7+b9IIpNb5NzfIgcppJpx31C48hugFnJvzezEEQ
YGrmKRmkLVfgny4jAyfYJTXYPAl7Zkq58ugUEhhHktzxjxS7wU6LMJ+LEWhU+ff2Xwf+TsUg5Xdf
XqAjMIUwwYRZNAkUXuahtEpaX6LksCdf7gq0p1nLfO3WqSc6W6l7RE1qkU4+eybX036mDvsmBS6n
WnxcSRwJxAthPMxuilVF5Ke5qqA25quLbIay6CfCsF3aJtBWNMqvLPQ+yaFeWG0D6XFFgwKAL277
P1zXw5SB1nqEyreMjexCO5WzMyPbRDBGAT35TLMYwMtUOAgRiNNF+zlg1k7FwuEBIsRg52hAyZBb
zcC1yHD43nyifm4VV82SPSrpQhBhvYmeBsV+2R3ds4as7d5B59BsZ4wm/6W/KS3zmfl8kl6L+pIM
BzPLhQQ7E11+DyXjB/6JLVqoyNi96UDEBn+G8CPFvt7OFUAAIHy9mW/dDRDzLf4GnHHrnSDLFxCR
UE/1evQ/ho0HTu2bCx0ScXv0Ipcv1NvvCyoGbxVio7G7Pe9U+d3DJtl4GFN9mgmwPcIZt0XZpCVy
s7eNuVdvgApUeDliZvkO6TT+qE4KE0t2B7WcGIh2KS9UVxNI9TsPr0IfPkCnujYes0xPrBIz4wyt
xMa8MY/eqPkPv1Z/5879xcUAZYrkYFi12/9g1UFp3yhqG8HC1RKLKOPQ3z6roY5kaoLKItjpBxl5
uE9K9+fBBpjIWZMtskH8Qd+yfx4oIEeh+PBOyVlMQ7L8oPWCPaEc8DbMpA7RGOTg0yNrLncruTNx
A2H0kgjL8tJEschrnXHzg6hkqf8x8Dd41ZdeHNQOPyR5txHJ6XCeBjZTC0m014pLogk6mddjJ/ik
K+oDa6Nq16AMVe0QJzihVVrXoyUJ74QRBwhkcVH6k74wnWao8IUXznbwEh/St3XDB278CzB7YYm5
X5VeS1uC2o6k8bt+WCPW7n+1egK+Url4KSlvjVKRbkhzXZ4bExAsr8hcd9Qdxh0sD2cYjHYkb6jM
1HHJvs4EXNjukfg1q+xMyse+pHIJQshw0QpQ4jkobQtnqKaQ8KCgiR9zaWS7QW3GjawSjs6jBFZB
1WCzQPmkY+JkunSDLRra+Cmycf2rKnDDFzGDOysXYJw7OyeHreey7GUFqaLewb7qmCU9HuhKzfWI
H+mOtw6igdEjkD5a0YSeMn2EZR1EkaYNxax6aobgSCDDsdwM4sbKgX6d43lhoSo+aG+GGpQTu/hN
Qww0dIOIxMIxl1LAo5KzXtyOy2fi2yme9tCIu9MRjIHpiREc/SitaiUnaTOrXsJSIdqB/4biXmTv
xlKXuVALEUA5eXztoKKxCkJ93xj9J1eycScMeP0Fpq7CO5mruu9hIrLvk/HtbBRxFttQXBzlwbEM
87l/k7x/6Jeg4qjG23F0xwXv7dAUKSPru0e0M/aylAAerpd97xW8kNR238opHGmiCAzK3VS/7KVL
1RdK6t39VFfHGuQO2fMoIWogoj1yvWvYfEVyDgfRLFABUCxds2tqY56RPrPJwZSwRgtrETvwXhy/
GQdnaAbaqtpP6208wIrLMh3KPMdkVpTNH/1kz/cb2Z7yanIdx6UXOfuqoWKbkBhzdHGwjULIgw5D
tqnMVrATn22n4maDOAtajeyCWjBLSpYogKokKpgdaugAzteZg3kel4uy94kgyKH7nInELdOxT0NV
8LkF7qHRindduQlqX9bm8pQwBWDoRGArNyMFZBB2oyF5Dcnb1GAgo6bRUcf3TQtDydE3K2ngFgoc
cqefAPJEhVD/un1UpfmfPXl4hZlvrpN4S+HqMJRm1rXOgZBDYyofJvyX+MiMlcmNuo+NYmm9wXzY
PiTtpTV66seaZ7IeW9kH0bq9qlBgSQtr+YrhyDwsF6fLgh+c7Wi6kQXcfSg/GfUGEHyfs14UJW/A
+qSr/7zGX5JKrLzQiNhFikSKMfYcLynyM9zmEKWK0lpQnI9zzH362YEaghOFTY4APcWGnnCDUPjw
+eWeIZMobplZc3kUqt6kPhDB+T/7QuHreQGM9u1Z9iKnXMi86kDF1oN5G5dEBChsUSE5Xe6fC/PM
oiW81bkRBxjMa15FJMWb9fAbvYCzT73yBQvV9cN1orP3yGdhN2XB7njH2519njscXPyTmaS9dpbi
8xaiNSCBBZON8aWmu3E24pmGl0eYGvDLR42IWeMaDPhXpO9bidiMN2wmzx70iaSOH4tqjJZrD9Jl
0PfsdAREbI9vJJB4842anIKkDQ6OKxYpPPeU83vBPFTcuXZn48uH+mbP6Rh03GF+y+lqwesDC/08
E4v/EMobsuefgLpYvZwOmIH6tdnRsxM7ae7MBUrl40WHIa9mRHpuRhENo5dMeZLVoKYXoY4rMgkb
iyFF67Bp3zqwIf5YUV4LxmMkRY48U0FZkg+3/494MnJHrPojr3NvAL1R7GTiMhhTfp1UUybeD9jg
6ljQQKcc2BPzRsveb02GYoY/2Uo3+mPBQCxt/KxYr7sx81zMY9Wn5QAyHJGwul0LDiLOa0EEK/5X
sRvtWhEPQGTDyyO3/8dOcsP3ErtQwJhe93WRIsaWS1iLhhpXe4/4U0Dgz92KYUaDWkYvKkzlKTFT
2vk6e2apxx5Y4fcE8D2qyogkESQ1NycHQyNjAX+g29qHs7Mg7JA/jivS4p/lgKOK4atGLEqEEwtC
Jg1JWD3EoHzWt0lFiS6jxq79m2OkVSLRh9XCmsiAHqeRZonInoyEGAQAmrhQUWE2DXahyivENj2X
ppEONRq1nZNROGU1uxmgPn1PfHP8ZbA0IMw6sKAcr0vAabhjag6Rfw4Cwl0dPE4qCFoUpZUk/Szc
oH8OkAHXR7hMKS1Gznf/G/BWw0uJFRXJBjmqWUv6yGd3F0EWRZ18G6+XThEfmsJ6qM7hJ8xoDCtT
CM1C7smCf/IRv/xzaN9BhZwLTp/BmR3SAQBAB34+bLWpNZikjYHgBLfe8Ee0Qr8YPQJ+05Tym8CG
pZswyNzAEtTGJpeteB3E1ED5JRA/c1hk3p6vIydcuJbieu7MdeYl/SSoGe1CHCFdnQFEVFeG3oHI
QqbGCpPGDLBHBW7drFZ7w1xlJesbWAa1mHhdiWG1ZIhZBZ5RBni6X7/9+iisO95caFebCe1UeT8x
+rf+wMbShXxGnldL9piMlw7qTIqsJ7nPJ0li82T+xUD+Aq/hQuugMm5dL0WpC1zh6b6Db4sQbYDP
tVK0DX/MF+e12266jDMVbGxbYjZTdyYhIcKC7d29+BNmaS8fgXqjYkgr8Y1dvmCqiIQupi4bN7FV
Mdw9Z9IbJi6OcG1Vq73OWOEA0IM/nhf12WgirDlB3FIvD3ccHLREDO53VZyKwrrmERY7bC9BhR6c
V8CLEzzQibbO1psERtXQPONmZUR2m4bUsFn4FOhMV0J8880N5EYcpVheC5EKbYPc6DRNiwrlbc/f
GG5qN8ovrAf6GUWvfFHyzQ9tshtXtYQ9tZqG1zSOcIX56WAK/+1m+je9eVTJHlRmDrFEL8yGdBxj
8rXvF0opLum//P6zHXomAIJTPdy0/9dVwIuh0Gz+wns2EhK2A+chtz5WcCPbCgb1UDu0Fb1qn8as
1hQBcfJoZbGC4j8pENZ+iu0FI481LlP5Aez100dQWXFd7kIgzoneoyEqR6t223j7ToeIdfOZfB8l
/OqXKSKMVvBddautGDKg2gqhPLAFcCz05myQwk5oxp6m47FjlzhmZVNqcBkb67pBOfG+6IGM80Xy
LXWkgeb5WZHoSTmO/TaEeFBPP/VhzHWehxziPQ4+etYT5dT+Uitjg/s+ZHjn2I5X6D3TzDNposl0
U6PrQTx/oZd7KRZv53mG03FkfbDBFYIxA8rceY8bd4PIKQhBi8iXUPXfGlIyREJDjZd1IItHIJ9c
oOjZ0XLsm+RQ4WqfEnm+R4EBbpnWGCUChL2SWKqKfxpUSq0BhxcjipbxBy7kPiebZQvZ0MvwLmNu
Q91biPHoO34A3Vbi2d3uGTI97ju9eUnhcU4Pt//Q2JVG9vtRasjxbSVKhftf092UMo8UBB2v0pzo
J111O/cg8/to+ojvS0wf5GWTPBnCXcE2TzGkJQ5og3uMNo8P0NPVvvu5cTxm/Vy+13ikJlQ13xoF
qtv5s8kCfyC/03sZ2qGZSf07oaPkAqTUOGfX4cHAVixIymxZsqjW/4usjxkG60Fratbma4+Bh3OZ
9tvx8jxJ1wUR5/lQ5U7Uk9u3kR+zW4U1c0OSTatOLGJ29xz6OJkhbaG+lJjVMb/lQM6km/LzBlW2
kJ+snJDAwqFl0lFHef3Y6jg71ikWWuHd+ZPCkT8V92bLoqmCgbV4EgcC+XeLvilwgbpGmEQ9x1AB
oCOfqCnm3OsfvrnQKrsnoLJv1JpjpS2fxkyeE1+a6/ayEXA+kRTWkl/reOyEeUluzyBeHSiTH3Ha
8fBp56lD7tBpjWOdZ4SZzNFKe46CLn1S6kTgXZd8rcLxFlnrthC/NVj7EcX0ocSxHYsnpMVTO1/d
aqR1J7ppupXtUOUeshTwBF73erfK/vT7S5OeeeX/NbFT8oFdyyiZX6bEC/nFGPhSl0RBSsY/ajwY
Eudse1bmNj7Go2/c4OR7rKUV5wYUxAwhtpGDK/68D51MRarGOdr9YrMcoZH1w0ChYngMqm5aVSc4
JyoshHL13e39a0cbqHpndk4PMCeUy9sfYZN4zri8KoYNNMjC8X3VgRb+s4vFeKTcTJbJfqv4Qgtm
Rj/evyuLkfhyMRw7GTWG24XfF1p9vgiKY0hIf9qp3W83KO/ApZQMmUymvYJp5v78+Fj4UNeQ5vnK
zMUZ0//sQE/GE5QhHR4L6vEE3kRUl3nB0b7uSJPteg6x39Gq61HQtF8u3rnmAlMLqI076of7B6Jp
yEhtGT/sCMH0KAFY8pEaVy6XLldiCS4iqb5rgWLlu0bmM/4MrOOa+dedF4B8+WpzOh12mVlmeTLi
WH50jU6MpyB1Ix2weji++sUPdfzfna9/XWXH6XCKl8VtiFicM5mZ0zHnnMcEt3MXk5PNTYH1MImO
J00YPgo2dTEdARQcXX6tRZM8hh7oEYssnZfZD143KJjt32JatPTTeWNEEwbmcBHk7Y/qx7ujtqru
VkXMWdVoNb5nnJ/Bxv0D+HOYftitsHPx+ZcYP+hDinnmnWjEk5xF/u2C1lugoRazWu0jDYR6rfQf
DnNH1wbVXjNXbfBHfGqoivwDvoYxE2ibyPWW+qHSTpJu2ueeA7D/1J6qOrqZoNJ6hPQO1kS6f2tw
2tORoOpz1aZveAyGbDiimpnuRNvzTwMhPtZqxyliq0AmC2dK0RPRQcSgSBd2FWepM/HnopAINLMe
cEpJ6UBaUVz8G8R6SiqdzX+x+lGqxbbpQH2LWnHdQOW0h1DxBgsYYCZKxRekKOYJ7iW2vwBw31SW
ZYhQRjXlOF+GxlHtYNHXFiVtmLuQVMLzf/IqZ9XK0Ry2C6n7d0PNDX56drHy0dJDO0y5L2H2hgQ6
M4LpnyL3fp2V9JfDZrh8JBWF93R96C47gChoI7sp0P0aToiKTqo7ShLmwecxqw66HVlOJ25N7oXO
dy7DNnk6njRuAETQswYk61k2JddAz1mwx4TSRN837NQYQ6pKPWJ+1HwEV6c9wrLSCI1NrsXIT1T4
eBueATusyUX3oK1USJitlMG21+zxJmN2GGaHy/EVEOj9hEw4GHdGhZkCZGi6RAtPkxGs44v1IQWy
3Gd4kukFoVz4dSayQ6QwK30XLOiLjiJKpPXkO8KirY5mV44UeBPvCBqDb7MTgzi2olJH+oSoFmL2
CKBCHfxQDHTgLuBgLktoIofo3bO6Z4Vkd0T2NQ5moCxv2ci0X4sROXTeipHuJOz7LJIySt8H1PVc
LQl74UXz8QvgpgezilQhqRzA7Ea4jPzrQxEseO2lnakTsxiTGNXmhVL0o0D8Ri17pbnLq874TZM3
eRxbUhU216sEzoJrZO4WLYDjoGrjb3XgnZUPYJ1/TvqHjWHs6N41XN5R0K3EQAALZ1QYtQFnoxkv
XCEeyeesYsHLtEHdqIehxxaOiMB91Osgp8EGbADmquHhJMO3sb7QnE1k0rZTyEZQuWoPkmy4evia
E0KMdddlQRrr0bxVHHwjvc2xVTSZ9QLl2/u3ENH9Q07gJ8YsxXVgM+QZ3QHz2N1QvWbaipIDT8g/
Vb0+j1yk6u2nRv+ay5rG7/cOulRb1Q+r/w9tDVDW5oZpXrlkCdgw8C8dfgi3fP8OSJU++eFEVZTb
kQuI15Q0I+gOHwFxLhzc0igA0XIGekeZTSNBuZ2uV6zZGjm1uZ/kOnl0L4E11fxmR/uXO3Eosxf9
UmZ+bKMURtTEJcmsetMQLhHWhsYAav/Qrb/+kCs7aUTmPygmbey3WgPzjOh+Aj1R7BOjvOw3xigK
xpMMJHfzluwj38rNZCSqYjOzAeaJelZJY25luTgmk8I1tAT5dM7ZG2BLTdBJEB0JdfhqeU3+kejv
zlIaQStVaYNwZtFgT5fNAbfIyAA0z7Qx5v24qMHptHk31IR8O76pRXYJCSmttQonOF9REoBty5m6
DkgYEt6Cg3ZxEeHHgT3xeCSb9aDzlAgiqnEiqxqK9Y3SgoZS+ym/NFRs53LvjDVaFxeC/o6EnMll
yQxFqLotfdOZLqqRBwzC9/XprBlYA3zo/RJLzrVCc2VbIk+RFiTvzu1DMjaiLov5F8d8fKbB2ypn
tAoCZ4Z97q+86VHs8IwoAd3GRe+hX481FRjGxQ4d74rMnJlZEDlKmeCEXp+5vyIAA5Uybdvcn15x
N/hms4PITpMOpzNLv6zn89uKfuuRDhf8KEt21G/fAJIaedjtMbI42a4eoT04SHpZ45E/4LRwmHB9
7rR0/1qmP2aEtx1m6+oED0+dOewHPAag28y24Uaio3NeeiOGDCLAUu+VwnA+Ja2pF9VaHIOhEFXP
Bik+MqHzPUjfoADgJF9Rjn6/9v57wCBZJ0m1roQaDcUSWEfKyrNtMwKKNOHipTid6h4FFObl8XQu
NajxZ7Peg58svQ4z+UnctarnJlxAvKk56/rPcyL1jIDRdD6AzN2ftV8IvanCROLsBonYO9N/AN/9
GmLldRigPrdX3+9pFsjxWkN8DIUvczkX8Abvtm21OIm+wZbessIGtoN940PfCZBn15loP2qAqY0f
yAEsUb3W3h87yxf/SNY9s+ZWTk0LWw/Q77ia/uCDHtzhwgXMsYld7NqMjbIh3njDgwr6sbg/FnCI
HxK5TM4SVNHchTDTTzNRy1szc+HpBr6BFZublGm7zFFVlSmVcoEQyhLF4kPPGY1NvQ0lmjRdM0rF
gVK1fWae0/vNRyjQKlqUse13Epd4aMRuBMugguj4+FnPELd/fZ45lKsx6+CoErcX5tUWNKrXLoXo
hSyeACwnrlbjA1ILNAY5rpwdZAogCtuWwMZ203qJQMq7xbeQb+kS8GRbbgFyqrC4aHgAQS9+Lz1v
iX7ak3UUokrrYJvnHAI47Rvl9cq3BpPC8YhjxQ6u/6tcZ0u3BiMkSReGNidFYaisOV+Iaykb2rQj
SXADaEtV9J+s+JajpxSIP0SI5F83OIAy1dNyMhwGIn4dfKrJ7rCnk5SJTS+YLMcWxmobU7q6twGd
UopugHAajZdJhGh9X2OVjuyYFful3ZqF1xgNktX8GDjYQT7rT/63pfXemM99hTf+ImC8/HseakcY
cdV0djS1kGJOr1xOElW73vfr7mtFTKw1g/rF78JXIjLP3Gm5hJvX6L28DZF0xfqzBoD9YNdtnH1g
Yd/6qRL/V01CgQbe8AbAo4YeXBPkIWLj5FoQlZnSc78epr2K55E6rKELHg2kwfpQlDxclyqtj4A9
lwfF1cRn8BFjrt7TiCOKarf2LXrDlHQeCpHbzGBvtwldf2JzJjTOsvBLzVT6w41xtbJiH0etj9YD
5R1BZU90hAA6M8QuHG5Lj6n8wTmNxm2X91dnzSAPKvNtlNnqI9Dai0WuUiHtzCQWw0Bia/UGdxhI
Oo/ZJTig8Rk5UOmBTNEg1PoGvWijU3AltBmTRkslWHxc11iHThx460/f0TSdUeMeAPaAAHk52RTg
svAtjOtBcf3ieNyxs0PoRQMtvGelkGZTrVZeVbIJKLek00rScJ/ZBuzvPnD5ikyUp9TjqL8j+Aui
ktT+Q7an2ZwSfFr3zKympkvK5dBY/3wGkf8i3Gict2B6PgIc0pP9l1ik1HtZB1W46dxQX97hejJF
YIzcJOsC0+/QvDF+v8R7UE4sLJ3TxRukhhKfHbH1vfFRId2IW5KX/V1L89PBU3jvs4MwJxcnPhQa
os3+sCsleAou+ciCL1MV+PVq2J0tCa3f+qGMQ5mFRGn/bvwjGvJEqPG6xXO6rEb5Cz0JNjihsZTe
k7izPMB6xN29xXrtLIr39C6PYbCAwtrUZs4NAgR8M5BmhBSqBvqMY/lGvJ2xbecm9mU89cKEK3u4
PgMIC+o4f22cGD0FKH1x8G2MdkIiQKB4n+iWhwM67PHaQrChY4r/YXlgj1LDCEZuTBNMV7vMujRo
InxYYZ2DhBzQCrx51NHs/yxTe2OYrtWJpcYO8I1jrii9u2svLXEl+m3LPWUrVmG7J1kk4x5f/scL
XEkNolQKApmN/jhCEa0YvzX0ikRwVv4gE4RFBvzREiY1Q/9UjXVG1+A8i2a8D4PPjH8DCnwIk7IF
DKsEBF0zxskIU9sFPYqottnsGijBmviEgfl1eJj94UMFTCYS5LcEO43nWiZJmmdquRcLMhNo0x2l
HYdTFzfjgZs9hfa6Vqaf3vTXYIzulYxYiYzo5UFbZZemNvOfnKSdX+QP2U5UJ1657LwHLCPfLJoo
runBpN/Nb/kMH8La6Ku6gsSzlD2GYEY5300m83llnF1Vookbb/arxu5zgiu++XqRHBvnu37nQHuR
Tob4D21+hHNGt1F21eJx6ddo5DcyqfVr6SZSC+uLi2soy/CuORtDA4/k0Qb+dByFcIfhMEDLYZP+
zeylEJC5B5EtbcRxB2/GrJknJc7gKlK+moxMAN/RfjFoxVuXudQcvqzaTi399livDRO6SM9Q/gAv
0xWL6sYN0V5SAS5dZzsm8H6ZvMhIZ/cqP5A94wRnngO8BltiH4cgmQK9/clX0ky5SCnsN39SNJmO
0vN6qYGoFAxDxao0eZsddxZzGhxhZLPDkspFLzHIUeKZdsNQXGgkRfP88XxZivVg8TUCIvUbTZoa
luihum0nuo/LPyelUy43KCM/GYLlXOZWvAUStoKfxvr2t3cJKADyTreyDOszWHaspdvJkC75+ls5
deGxzbzyktuK5mQR3mpNx3hMXohkqOHrzQrzKRm+OHWOScs6dOCuFIgNId7/bSswsuYlGnbl0h6c
5IEIonwviQZmoQAE3iEULGBtfb5Dc89KmF1yWkeTq/+zr9LUBHz5oFKZTho2n6Z0DUhqTlIkWhqH
TQLUbOOhTErlI/Qu5X4ELUJUFxGUsgwikm8zC8NTIUCNEC1lPzheEGc/der/IdN7GeTNvgNzDV6U
AtefAILhoDK3Z1wXzLyeam55FGwpkysgnz2zs5f7Py3d0qQ5upeAzMZg5xyBVY8fRcZrfcszqav0
G81ucVB9wsb1VHwk78m3dJd0JYYi440+pBCiH1pdAZ/hyvJkMq7TKe8UIeg57DUZlrq+oURJX6Un
ZCpRs5TyUAtAg23MbBASQFBd1/nbYtkCA5ItWbk9Taqw7Oo3wROd06eSefd3dxhnGlbGf7b/HeWO
Ahd1XuC0lTIKLPqHGFDOTIGu8AC9dw8uk3kgaNctHmztpi7/0mSCkJSNNgKWzhD8Rj9Sknpbo4m+
oQtuJVnSDPix0JtlfdgTc852nucwDZTQg64ITYFOlNFi5csbiZ2sH7pT0V6UFT4LobedsF5AQN/n
8JvefaujYNLM2vU9wa027h/GdQEx1q2pbkM59sI8cTMoj1rD5jP7zOVBCKz0NqzP98UxIcMzlEoy
JLcymcdC+VDhQy/rGJct7qHOdZWRKh4B/OrafcoLS7OSjNx8a3hvFwOW/nYf6Iojj8Q7wCeEGDY2
swEPP1eSK9ePGz17OKOfCnxQgtKvtEkVnIwgg3XH8Yx2NRBVis8IZCKxxJKVv4f/N3irsEiybPbs
H9OIi0Wg2LeWT9TLaLdTWyp6u12suzDc+djBLj/yLCk1go0E68e/dSd5NlNrYCi7avz7EjsouHf6
tQOdt39Sqx0j+YJIrBP/lYAnjMUv95BTK1RlH6BPM7nq3oxyIdChS4Q97KsNuZh4ZOucI5oZSB3Y
tchA4f3OnxanGA1YMSkHmLdM8Ih7ca0jwWIiMJSXtAOAyclNDgP0o4kjWabir9bi5l4xx3aT2fJk
oRValxCBS00AQwIaA1zEoU2olZu0/pNn/GhmIQPXg3aH8Ii0lr/YI7pNkDFFTslfsKQTFiWe04qN
6WEWg+QrnL7st5XGAtyYa0VJwT4HyHZihxRKKyKGC+UQE5gXM8Nn3i4n+dZLzDpkV1p4F1jdwNom
iaxSqply3zdq2M1HF52zJlvKj6nrA6c5LPx2esbixiv5JAqyQVyyPQGgFLCH8ABCj5gcnFcF1Scq
sLNRFfri5QSWB76gbfOi4ze2HI7kh8uWwv6893Yp7qBVQsFVMyKvxk1X2P8zU9C63ShX3ePv+hY7
kXhjqrdH8vDomnSJH+PhTJpQTDAdJ5GSV2X0+T221eFF4OecA//SqR/lYrJ4cTemL6/KuLLlIGI3
1RyjCf5CZ6+RXaxi9qCP6FwQ8jdmFG4aQP9AymVp3EwP4PAhAzFqJwYJTIreiCvKxptK6rlsFsWr
TF+YKLF0LpKQPLjSIt6ZsxUGyeeso2R83lLenGwi+Gv4QvtKYc4d2YGwDZTIXs6GDuSPJQbyhPnv
J4O6MiMmHrKNQ35XVetv2WEfLPqVowFY6Vn/AGcY20cT37GHUV0164zp3mAZuS6NkHVmQfHoNogu
jy5oqcDzAVKDcvFhBbgSN7++4uo4r0Ct/6jPTTLF27WslTtmjvRdjxoyeTp9AgG+hXnpNQgX/rMx
CN4fW71qoVdKYcGhRDoDdj9Ey70gHnOz9IUTWrIDbg8RPcFgmjE66dgXkL18tGr7qWoupSTQNBA7
X3ghDOMEnWRZ9kbUu4Cp/veetmfmJTu7szRIkNvFENnCtO9+AdhXH6qenbrXs7R9ffKXavA6qV5X
hyvXZUOquc+T/IJNYD2iszN13hJ5HoFhIYFbQV64u4gkWC8rqpSdM5TAY7dj+uYQjtc9IfpO0/P0
kxINxwPmnTLY0pOY41nCQVxgxPUgNVgmO/ZGZO0zt6c8ahl1cuts5RyoA8/qh8jQF/Xd/moF3h2v
WQqvCv9yiTeSVR3V64m9Wqa7C/vWzC/RvL+GWPcUlAA+zNUUw/hqsdbY6rkEpBrIIbXZnXMN2dr/
/OgOGkE2lE9Tstuvvoxv11j4Ce1QzcgLanQU11IeeG4j8bEs7ILIIgE1KNF7vHmHYRY72KBoTjDi
OQLO4MiJFhHuIyooBocQuU0mmTXLFTjFxUEGWWpkDOWO1oeS/FOmddsvK8zpg8Nyqy/taCUe+ACO
B5TGAahleIikV3iFatXNtrVUQ/Z3lyyH7Y2tUYFerdHBKskQr/2/fUbEzNnC5jBRJERdkGBB6b/U
koO5rd53JVa3Ib0+X8xAdlYCIhKPqUe2tKsCl3wDQ3cI1x9477i0ZGpzaASF4runKSHR1S50Kh7W
ft0AShDNhSUw96q8VXayo8KVW6jA/2e25z0c+O+DzBlbq5lRr030HzpBxdpsRyXVjk6/KqoSNma9
7+IDW2FIJPuTEFNtGUttKF5B8/2F+UJKE4MszuM/vGQ9XaSpmcDnAhhPFZOadYKRFVmj9rO8lfu2
QwFfRRPdBq7HXsOmV06GnXcGF9dWTDcZn/G0B2WAzr+4AzHiNsI8b+tbBtFWtZ4TQRNcyu5HECO8
O/IsegwpXMgBKORteN2LG6kJbiA30rOVK8hvXHQC/4lzoBV0n620OXmje1I31rdYPEOHGDVojjwf
UinH7cH6FhyH/YhBd8u2yPCJ5rLa4l/QtffnFbFzEt5ghm9MOJ7PIYSdCMfYzLHOHMJc6jNU+khf
yQ7DD0vabqUCSsJXRddjskF1ZZAYl1GhmaHGkH/cVW5Fsma8BEfDlAkuCHXtALinlOFzfaEEQ7z3
hum0M2oBZ+lVbXIhC8R1dN4Oi7V+dltaqy+idCFEveP8kepwcy71eTXQp3lEnv9LYjCGDrIZakQW
cIPOGaMzBI+afUgrRJOEOLNGJLtzeGPMVGCxkNOtddlcvKhhIt8OSTqc34+5W4gBVtgfauH2Uy/6
cLgVjNS1wPtd7F4yQScO1xLUoc1Z3CT/c9Ky6G5zzugMh/5HO0Lei0dBi0T8liKJ/jS3Sd3uYeD7
/s45mW7v3YPdBSXkM3K+UveQkeymIlYFC86birLtNcgj0gWLcu65grapbZwXUoVzZdYNPAh3hnxp
nqHBpx+LETwuAzZD3hOZ+dX2aBq/PhrCPybIMYys11eaJCFXYAhunysHtWSrelUgd54dIgWEZb4s
1QQvqViOc5cK7g0Z9rZr3q1wa9zOxVCbjo8YxKozw3hAo7dB8v/5i4M4GBHWwEGfZpE44muf4nit
62yjPGLC30zJ2kXLaFuvOZ1bEx8kZTYfKeXyQLSNCwRfWUahczeNj/23O3LVvVoXoY1IdPtZb1XP
kOfqiYNCfc/m5v0Q3fOWv4ZdNZjIwBNflae4ECrntpC+VeLplRLnjHWdBrfcrf8X/oVMj1/CRv57
e1Xw8CFSBm/7xrH2ktKnhSyFlU864GyWl48MSK/dVHALffwSEFK4JCNmNoVQmdHmQucqGXgeh8YP
+Ymx6JJDs90Y/3vEN3o3n12Ljqd7hPb5CYTSReoKwD0K9tCEtogFuQPHeR+bt6RSZHL8Q0nK52f5
UsvgBXv5QrwNRdxAgLJEBg+AgDYcLPDDqmH42Y78TrMxhDcElvfdvRJsY/VrbWnSA7TAjc095R3n
yk/uS0oaosO0VEa15B8sVbesTf8vxkjdAA8QbR7DI75+2fpQOhTMK97yt9u7WCaGhZSVmtELTAws
64LwTM2JYS/mKuPqvp+YSzZ7CM9t36NiF8UHHrSR07oTLr5fjx4YZxs4XD5l6SjuvAr45Cm1AkHH
TysSSZoP630K3rawVUbBj1WKg6BNVQTjxvPRJnjRt7gT/AEx88uc6RjWLVVPq/YhHQ+L9OsN/Top
uJZEu5ai7kssxSNfmyw7SSqbbQLhGUXH8atXuNWvtq7q+/jIjCyyuAdJsP6Te7INbxSKMVFt8Ytu
cuSZDN1Sxlo8lD1Vxlj6JXi3lO3YxCzi6AHSvHbpwY5+8LLNyhT00tmEs9T1L69Vj7sFCevyUIPH
23cuxY6IT4Z0Ubqkcgugn+1gy5KNsKXrvzNcOeyCqlYg+RIS+N8mCKrTUR+6qXF8aGdTmpufMHH2
07sCSMqqeGHRxQ3y/55C6dLduh5UhLaenTGuhyNSP2pLzh4hzFB19rgxkxb1bk+lH8reZbXUBbDB
cc0Fhtvj9TiIs3Zr7mmgAxKx87xxn4w5f+0OKQLfPaAGjRO0BFosgL+Jqfu9alZr40rdGRyRTuyN
xwdDu4XNlqYY1Z5F92EL0KcM26P37kgiluPTUZNeyoRL3FOyBPxjXmV/BG9vdxZ5TXR4vRCP4l9O
OMPBCEUBu2agPz1qQZmc7jnFZMhTPmY/coxa1wetb/bYajFyFJpCpljgR6NqysjMRpj/HQbYvV1Q
Bcr7rkpABjarMXuu1RGWKXOyyZugGix7f+82JJ65Xy9eMOvCzXeddCSP49Www8NZepFTHU7W5CTW
eQs+Ao4IDKAGkEIy0TKlApoJWl0sOP6mhN4LQ0QMe07vLoe5pltlqCxpM0ytZZwcDcfpo/OvQGmA
qCnhJsoHjgDKkMadD9pboJa8W5LaYMkAB3Hk9OiHgWueCgQ2yzanlmH2xyLejaioclkcxyq9wCiW
hX5c1v7aIwIXa9b9ihxDhKLsMbDNNGg+GkvYOpDGu9bDry+e+M8a41dVG0Dfv+bmaKAFRKwJEcBZ
orLUpt25hKIYxwno6Av1KiziWWgrvJFeKCD0mA2BPLqnZYPF6kRgcnxL+I8Ij3ZhyIKKYPDil6oS
nvj30NWbGEqa+LbFs8E8a8JDkWg73D9poCf+5x5v1JLXYbDuQB02gswjP97p359AC8Dr4GHwvgND
kVeHfIeZwfUfSFeG6Pv+CFFc3B1eT9fikpw1ygSX+cNV8zWRcMKMo4b/+TvOHIThMxl5LWFbyukI
FqQivyhyCZ9IZjNtRIxQBMdUnznKYh4JePTZoUqssr3YgRctGfGQC5UFK0wfYSCjUp37qx4PC3oE
dhMMAsEuI5k0Rms1FxofFZG214oVrM3Uxz29qVL5tvVGE7GsoXtUNNChIWfQy6MwdvnVUxdjEvlJ
jXJ9yKAxQq1iDi8fGTViuHMw3gxWUi4rjJ2zsuOzt7lkdVcyH+mC0syCRXXAwFi7XUcCKllK/+S4
hNXvJdm0mQrZ+0uGorES3aB+3J50HFf/PqKfRqyxNZQnbZ7FJkm9ZLLgfHerMTnjrBbeSCAVLQgQ
/LVHy43ZwimTJ31Q/W9D7i0Res5oeBpEyMA6gOSwutsqtGcl8u549u48E5xngnYF0k6WxR+q/OQU
BX/5hEEkP6zBZ7pi7h6Aqstd94bECowGAM1gApzUlPi4BluBeneyK8uAmzKcVBfwlrOhDEbbskuD
nBUbT6zt7wtgtLZVt00k1F5AB3/pTexjEYZEycAAE3tAqEJLvRuOJ57llTiMH89jmX1AtyutZq61
EHiqeIAxcOcqhVWOCCZJIyjqheFe7ECxyLuqatM7vo+qSQBKJ3aDbT5Ab/r3OO41syU2ILmrT8e+
AuPEZhdn5y+OdnSYaER9CYOo3mVPhT1abPuALHasiVB2Z41O4+LsN6CwtrGDcv9POeB7bD4yPA15
1kyLiMFTLQEDVw9XXQls9lkouywySaWFz9Oe0TI7530XOFKgDwiDVWA0QQrsuQxDp4qLl0CqAsAW
OvR3ltwrJo3RKS4/2OH7MXsq4LRDfonRElldNLRtVf+4YoOE8V/En0z+f6FyZD9Jqj8ww+IHr3xM
SvQ/q2gjwlR+jiRh2+eYhiScDlsxw+BymyZVQ+84B8IgdyTO8WOfVDwpG+8J+DKV54g2tHZezart
K+0I9gIUaIw4PQzm4vka/7aG//MG3ZXxaDOWEq3SYLWkUCOXXuK+whMbGZ9TxgwbGxicWG6jcCN7
7L2SnbnK0R4z3bHstbwKLTAMfDJGmDpQakNUKFkyvxdkD8VdjwLgEUtHi4WXQ1O0O/f9Ulwknghz
adfEBx5wNHURdzjuxpb1zVEmdY0Mudzsy7Lobrsosrvt87PDYXQj5ZYQK17e33BtnOQXBgLi/LZ/
+vobCEdnLvjnWFe8g3z/yxd3bPoIXDeyBsC5wC5vB9pqI+3zHR7WPV1Efz9NKdZFuc6iZcGkffvj
kHOAq8IDBtNcHQ0X3ceMgKkBE9CQqy7UNg8RLm6hwC3Y3iw3Xh07ZRj7zUSUQzhhNHwF+7JhAvI7
m5PqwBM4ZayukZSqrt2lgUKNAzSkBRlB837nCem0S7L90Rq4xQMwVggp0EAcXvKVKaYEUq6w8ZKR
U0qFg+DLPlM17cUPkuEQgQyBdnoEZ8vPgBwNMRxWtKA4i6ib3OOmowAxvEGO0OK8QRo4s17wXM3X
twOHbSlNGGA3YYXEYTD6nzIciqh7MI2AYDpSx97811x4PYgfwuAdQldHfR3OZtNIXJ3ftk3igrN3
15DRc1oJ07FutWVP3Ro9GkSTclWLCbBWnqwfBEIf5uNahM0hlQPXJBjfRZYomi0k6CXajLX4k8lK
gNnMSJJpjVCdkNfy2XPCoIEZjuKA9HBRNw2V99Oqw0L47axkIFeK7DytDvg1TLAtx6j+5ZSACf+b
IaE1Hg2HPmqyxNYbimDGHaVSREYu3GRzikDpVD0gSch5DQD02taNoSqgdIbTrg1mli70cYqkohGx
LIbeHRs6X59cDVt0u8KU8Zh4S90PViCXRUQ9rL8PqmjNkRaJMgLHKJqHv36t+G49embx/btkT7Ur
9rrkyIc7V5Mn77b2ndcrMGJ+2H9k9y/CN4DKMH6Aac1lsCdiNAEgfgFeTsDwuHI1XaV8BoE9aVvr
sC7RixxCQIAGZ2F8HD/JCQfqf9UQh6Dpr6JHreUyk2VXoECqAA4EMlF+PF0N5/hEpTuGtPdnidDx
JqE7j+N79g2J+vs1OjWtQtRgGFFaPmRcUSEDH9nZE0COeFbk1CwAavXfsvUiVRhvLWtTyjjvN9lw
+FnOC4KBvEiHUTNyQzwrNpPpsQc5L0yUJfXEAKF9Lvx9t90uSGIur/KwMCN3Wx4WuwfHwnAZZD22
tpEncOtqFVT2FLkCOR48bK/tWVzsnG+Hy+ILlLm1hxSt7FVejScb9xe+vPXcMofsgQwStpWTeWZw
sJEDKUzFYN7bh3dntT/6F27EEW6Sj7+BfYLwTVSjQ/2uUeoNBYKZpVMhZQDQgSzV0HuiOTBjtvKh
rbl7pC7bHNQ4nvqG/qOpAkX2Td5oaJsCKXbqODYRopfbroRIry5ziG5zjT/jGZ2kSNgvc60d0HJW
TRtK/sANNM8cq/JWYUe5uZSG91tk5Ou1bseJV6ld2uElPBSezlSGpKcxbRtXGeaq53CJgEiz2CHm
WUwk0s+aW6QkdIrQ5MJbpZo0NNx6YRDYDg3k9gULckejfVjLl8odKzWG0KeUsDyIhPp0OeRIQIt+
a/UWTf4ROp3jWAs0ScG1RGpBd4wFUgZHmYyREFXnXlonWquj8Auc50XLxeSpYav/amoj5x+gDguj
+5jRUJeenhDPm59LuGGqz57Oz6x9yrY1XWjLlnXJnaowH6aqdCD5zGqMtg1LQWihevYWYvJGfArS
epJ6C/P4arxidFVwOwvev/4AjkMSWUV+QY0zFFpoU0BlRiKRQUWpKoaxcXfjgJEw4wHSM2z2GFhe
VJaTLbyVP7s2bsqhF6MzvU2/6ATiT2AskzUXtm2J7axo1jqVbKapG5ZbyfNbKgfJnzS3BNqMHYFn
biCYnRuiV5WN2v2nFFjpelxHj36E0lOM5WXjH1UYYdcse1PemxVB5h4pWy2umoashxVhBcVb7Y+u
YbVMjcdKiCAeCRc5ISOOinmACY56uUSp2vs0JDkIaKT5MY4+Ph1khjIjU8Fgme4D7oG7Edgc6zte
aRVxAhD0drSlMRB+4Fgwmw/t+UKjq+sN9yhtwppZf77FM5gUDLZMscLofKQ5vBPMN+y+17Dl24DS
xmfjvB0HEmp8decnpjr6O48ccTLzDMbueRAJWsb5ImnCkx623MrQsVa5chQx+XUgvWtKGHgvAyxa
Lk+J//TpwEPwS/s+Ux/FCV2/WPpR/35HAKDEx6IRxTK+rVugggPf5taI5oeNxMvwYoVU/MTQ/VqZ
OlCW/yAbhtt6j8duonssMoGZWQv6kvVA1NzUEuGaky/oznSrMairTrGQz9RbbM60zIQ8j7FKXlEN
JV6Wa2LzIyvK3pLYAMlvJy35SxfiOKNmDb/UEcfSIkLORrYI4gHXvrAVgVCpax7rzhFoWogQKtlx
0qA+WM0bOFIX5d58GyGgnWYFLErNqR9SNEWeMKdHYpfjlSP/johCfjxKzLx75ESA50gZBQOI4QEu
jpJ7Gcxmwgpce8JV1d2V7pIrsoWbcet1kyCFPdBsl9RGm7/FlYzSA1VhxD0AiG9OMvLwM9aAFzbg
qUzPh+A9tzSAzTUMt04okaOqi0PmWU0VOJonXgs7m90uVkee/TRvVmEFWVZFv6w/DlygI7fUJFvU
CnNNg2UwJPoQJyyU/b/csBa0mxn/550piSu7OEeiWYMtGiO5ErOIHGu7N+4wvSypAa+LpKSqcxYb
iXyku+2VC2YBWntibd0k921sfI1DAbn03Hg9pM/xyt3KH4uxzpQdzn35GOsPRtux78BAWmxYKFLP
eEXTT5IHSVnSQ8IqU2wGa4GQWYxDfuL3TISCNUguUJCmw9Fo6Qnhg/b2nBE7QfBrDJowMOz0qtxI
EE1O1/SAbEBySur6FaJlg/5tfU2mMn74FDwBOkTLDYo0T9D/nSGBtn+hB49Fhy5Je8ZygAOx4fFS
Mr8xzQwaGPdrV8ZqGnUydSYVO4octSn+HFg2ClWwesHvlbPlG0UU4G5gVBIuaiuIWfsQ0R2d8ZIg
7Jz8zz9UI8CuXmESJ1D/gpleyQvxVvaYAYnGStF/vv62qy2twNNEp0ZiWfTdjuPiChD2FzV7RQdq
oQNFyqzzyn9VD9TgOiGfwQVcv8MFB96OJJzSAl3E8fge3THRVIZZMa1oPxxOG0/p3w6H0AkpTkkp
unf3mF8a/lEwATV5kKCNhhN653xxls2VwpDEoBdvagj+JFMHNxX8L3e1jlF3gnmYZKRLvMNsckYg
BuOQvDGuQeSnRsvuQMTJuCorSkNDPkRw0GKV9izcFp7NLaxL9Zg2Kuja7otrXED0Oke6Q8l8gCs5
kBcFY5Le3eWPNAB2tUZN+aMA1CV2E0Kn/iyaEzE9kuBcGWteTvHhQqWy8q6FQ+fD2qEexFn/6ho7
76P5TlZV/fkbVAnCaWSGibPmeNm3NwPlKolk18dnOpX2Jo+hif44gnV7PwYDyTh4gEGnywF0ho25
QpEgNE/5X4F183OLIccaSmOWYyMjBUYGVH9XjMJUGuIyG6reHXFkjSjNJIAbFvAj7kP44vE6ITXd
C7eB+eD+fyGWwqEJvTtt6d+pcuoTxgxkm6M6R/9vH3DRSxgZoHaD9uNvCKvQHfheVifhV78aK4MW
OmCoJYgW0OBfo9ravU3ToNkfLo9kCpMFTvVurXk6ITtpQBYUedD/UsEwTVS2BpnlluW4XScWPBB6
v6s3L803vZ5XDyDsjwc0qT03Rf5ls0HOsQvJkEP7eOyIOF5H7vogj6VXW5asktB41zbe+7P9Wep/
SnKxmGoi8B3lhn1iGo3DauOt6pad+wT2PCX3LA6dGbZ9DmT+8zp1tsuI70DIELaYR6g9qL0a5dE+
ZDY8lXx9s4jCpLdhTX6w4rEKTTxozIgg2vlkYv4Ijmuru+dBb9Y/6gtPVRqm+x2gtB4DQ0UsATrn
xaJYgPQdotVvyTIFYuWzvrAZVyilt70zvuW4e3KjicVNvR5d7MKmbBrXvzQUGg7FQs5wZ/O3s7r2
BD6Oe2iuBOQ7wMbZt8CmXYgbvfj0cusEBdL8YHTjj5s44k5G+PqOBZky845wHr5nR/a1VLarwOLd
DAX2WGtSWA5Zx4ojc+XgJJgPvuQlOgEQNpeWIrX4Lpfz5kVx1ox+CXlIxdCjJWiTSjH5jQ/+0uwQ
m1mvvG2Z7XOhv/PZlldcITo7uC8+BdgMf4aO3Bo7FdmRne2j+SASw5ZacWAdbZQ1fY+dAGMatvSv
p7Cm1T0ounXq14bUHIssKts71Yh/HK58zm/+GAHQ+4V4cLvr9/HfcsqyTF5kg3Bgq2xk6XHYs+Tv
nEB9TvDqjltv1OovVcmA187fAu3CSVc/VXVbzUu1fOclQFtpcABuNI00i3n7Pl+p54p8zRvpqrl/
ARjTeEIk7SrTl2VrkrG+c6MBLNrEVZJf3BUdXvFs52M6bng4Zt/rMKu/5O5nsYXkRRHScYcUIkR5
U8XrrSxvcfcZctweciriFnKJjBeGWrQZ3hRy+kuMB3YG3GCuZnoFxooKdVtOfUsx7FT9TEmkomw1
QpKSU1z3OtxuMM+y1HCjZ3sSm8e2lreDjwnZomv90VqJ8zciyWL0iph85pg2YjdppTZW4UkCpY0f
EneSyct+dE0r5r5+CgIW3FQcELWH59ITIuc4god2IiMxdlZ1ff9VwbkuOAayaTrlrnjnuPZqjhlF
BVLmEYmtAQyLQiIWHLaMLg3H2LApppcCE5Wa2C+yNsaqNxbZ8K9I8vXndfcXILNCEUMh3yvE3hX/
ikCeGa0Q+f3dFpyzLn6NfPSwNDS1tUEuMc0jEgTYKMepxQThlTkzqneaJtbQPNRVZOh1X/bGCyEy
h91wncqjHKvta2oimbEDL+fPYANv/spwc/e9v4ExqmqZi/slWXpkafgFxLoyKyDCyN2V1smBssZ4
UBfyC2Hg02pbHygEBBO3aLuhxuLdfl8Ym06AYNA3wgO66tKlzUCzPklIjnOOlLOP2MZBk+eooy5p
jE/e9oR7nDZc4v9sOHZritNxjrAO9diG20Vd6zM3Hy9L9Od6mo4HKGowDmZ/TExxNnPTKtHobKFw
40mkZQKwzVijnRgv48i+4HESNSpwmKrvzaP8UlS/KJ5AEC11JEDaqmTPzk+0Hk2+3nul6tCbDFr1
XoTu/PqzSAGpsqTjsrha4NgbBr8dw7PnCjpq8Yo5WESWcM3G8zURGnKfsLJh2pgTAu3KoB4/1SPr
D0ppyZq+5fdkk4coiDTKl9Tb8sa7aUKZHh/cIESHI2JQitCRkqLylOo1iMhsuhgXmexXURbS4tNC
ntO+3eI1pKjZFJFMVFzbd5CKPGAbjM9hvDtdvfVu8GoWNvi2S+5IFlr9sr8jzERSqorjMPgjmzCw
8xvBSRTVg/eZGILVujiEZXXej96EU789gkihiJ95W0DTlE0XUwW4ZAjlckoQL3Auf1wG5O4Brnju
6fPJgTIP4dZqZPlK1h0ZlAh+acwhE4PVbTQZUjSiotIcyNv7zWYvK8HA4SvshD99Im3gTZaqEgPA
l5nDx+Df2S95nprgDEWlj8mj/jA5Qa+KdsI+8E1TU1plsdWnUwztaliZGpHHbi+PjpgC4OMd9Kgj
XhXQjlvhpU3eg71uXV+vB/6FvS9VBCDjYGGNPoZKQsx7RAXu7OI4IS4DRiaZX3uNBLY0XTlCUJJG
WUqGPB1r8m98GUdC87eapP36/aVMoBsZtrDTuxqL5aV4K7uEyQmEgA8B/b4sYaoewBWFhkGOT/JY
kC37q7IDsXWZhEa02UmMtdMPGR2+cF/pA22K970UxvBUfMxjdKYhrPBzPV0kEG9xeDzrKcvjCLO7
gTXKtiPrY+9mhho3vz9Mcu/Qu1jKmbGPMD+/s3XVOiLV8YK4iquaaiKMyh4V9ShTxEf3nzPKKUBb
4O8Plqn35GfTcxnAIVFG9/jW/j4xnGgzr5+nqJFvW2rrj3j1XD0f9m6+9/3X85Fi4NbeBgNRJtrZ
URiUjhj+TjXaUjYSmSZRlZB5nKASy3wL5rIyeulZ+DhlU0X63Webb/PndOuFvuPI63LzH1sEHDqV
+4Bq4qbyBrWZ/9e5dTrMjyBJIa2ZZ1Ou0jEoIG4h1wm0GO5VpfaeLpx4mlXJkMqm1zTdpSDsJO14
9NnQgLIGnDVuh/cTvrsuSDePUSLwZfumfD7isYKKJjPfPfDg/xe+gr0asfC9Xo4mHH2fEAC59toq
JFHqJuy7WdMF34LuyIl2GVBBXMezD7btPvLuNlO/W3Vp2tvZxlNj4eoPrDa+JRVv0fFsREAA0uQ5
YfFNqZYfNxJCcbZ+lEAne0XO86XLd3h03fmi9EsOYqnVjuljbaRo8LeWExbo4ejiYH06q7UAD7SF
NxXa4BFytD+oe88Cc76gd2lr0yJZW3Q89pPa29nNjmtybVOJeXJyJYqDlpGweBnr2bgsWv+7Xgcj
Zzhv6JUGAN5sbrbePi2GCzUGyMbfNdTVLwPL7PkSezywGC7iWTjo/o6GRnOfCzneYgwvL1Wfm3pB
a28ZV6MYczgdvR4JDFfvNRGkhVHlGQkV/1XYfEsy8CeDcGeFe4tqBLMezP6aHpUVLx6RVumr8s8G
oiufNBP5x4Tl/Gg7jX2kWHOd5pK12O79NrUANId/CCdqYhEbaDjAGq4gvq+tjb0YlsSgC7a7uw5p
suHa22r4MUKoNthrbWnCICPZkL4Q14jwOWsZdT0NNB6XJb2sGLydolstLpFMwmfk1CHerGySIvti
5o2OqkhmlpQLQxUFpnlwdnM1tF8I8w4im74E78oRpt6pHKTQlDkMZ65kRGhwlbJ0UMR9SXy4/ryc
Vouu2/KPWySaYYu+l+slg1axJdQXTAlBnd/2YQj49sqXHd3UidayO/moaK8StAjzhwTzYyyBVgRR
gexBqN7rC6sEstMvg8OZBDniXcQKXVOCqCx0BrDRE889Q54G5JJcfPsklGcrikV/1sZONFG0yifE
JGFb1JsOmtKi2oVlKvjXbNDd3GAPm/dJMQ9BuiDL+i9Sv8A2as6dDAyaJc1HK2wcoa5PQc812q8l
vGOk1pdrS43K5vtxVO5rSYcMe8NHBrW7nPAfeGDpnhvKRvTqmcnfDZKuueoOV/X9LmdrjhN5nwnA
pI+7PnkozJYjx7TbX9BywF0i9FXGVZiaEnpLu4L89pRfzOUyz24W4s62BFGCalXB4SP2HRRMv2m0
DewrRCzik6H4BLHIaixq3OqI0ZI4p+AY05OEhKhFfItWORfQnQ9b6CLehmJszChRUVAwZIqyBf4P
MCOgfEpudGAID7sxmciVNCK/Vze43tURf6uHPT+UOLjEJeBgCUKyErYFBuLQ4c9q8gyBSj2REiyn
X9xkzAhYpHUWdv5BiGyv7321ODJt3VyDS2TPQ4d6awz1z4AdZhToCRiDqm/VQs/2gQniIs8G7YFj
M4XuiJfvLlkO3rVl/GxmO5aQMTn5KS/sBYu+Z1h50fxL36rj95LbUYanagzLbixjQvy57wyBwW3t
Hp0BDYjvkQTTtuEsozXhICb+sogTVrQcw5Z8oh7ta0Gg4ggilSu190nfIz2Vd3pc3xtP/IQAiNdd
YCT3b+9GmhnX+TsornpgCfV9P+7PDMjNL9nzfz05riRvVkc8xWd6FN/9CaGRZcGkSHE7pGvBJosV
vxX9B1/WfVr+jFt7QKMrKPuZHwx5K0n6xui2vSK/hGmugrzt+Nami3587Za/E0G1eZKPh5paWqOc
JHO97js/CH2U3XCEe7N+GU3cMSCgw31XwB9iM1IGoBtYEGu3xcd/mkd2mJwy6Ls1tO3wwgRjr+5M
hil13pAOdo6Em0vSKaQMz6ZlvgxBsDnXKXd5AliUEB+2YJsbkHjwE10H7vhW+JitZKZd4S6DAiEJ
LNwJdMXFQbUQqXisPPaQxW+2U4Nw3llcioG20TJz2rqr9JJgjdaYTdTVV7QravesanPUvlEsqsmG
rqbUNjQRD27C08Ye1IKRQPdUqAuO4+uiRQIQvCA4hWcFUTpedAGQtXo+/hy8bzkQEykVRdSxbOe+
exN9CSvTv3cVfGhbDHfO7fg05C2UQ3sMfpPmQMzR6ZPYMbXeXnmOoK7B0JBvZuj5R3+4a/tdEzp4
JM7zb0ar8zRSq+EXTweUkfvS+R4Y6zbewiR2QOZ95G/G8z+Q7ESZVJuI5/HesIjC3WaOsXXnMsOT
AJmkl/dxbDzBPiv03SaE39SUhi2usou6XLDnzp0lQzS9RrcRUGWUK+2iPZmLIz1V8A2IeVqM3e7f
Wu/gpLn5PX5dguZLbY7QqgovaDc7E8jaeklAv6KKjb2bbjnNaVdE86SBfssxvM0OF2LtLoOXrK8r
LCLvED/1V9MQQTP3jNbshFDONiVqwT48i5EpTHhTuRFrSpc67VeMeaQAdOWixIxuwVEskAmtpc4k
HHGucqn45w/BqOQZUxfvwppvRgp0rxHwLHfXZafSoMuMilsDXM0/gxI7I2DO8ZykC+MNc68b3UAr
yeButoDHtmfIq8GntXeo9TrxR4wblVwEkAfVePJ4Zix4kU8kwVX1n41smzzYFZwf+t/CInfAxBPW
D3kbzofLIrVsqZ/qHM3gicIz+7yW68EVBPxa8ymm0htPnnLrE6UAI/t6PqCxuqmV7I1csmoFTRkO
ydpLCdEOfnEiL9hSa8EJxx+ZVV5bOHTNYTBAAytrJW+JJFboaUgiPso1zSVGuf9X4tyQKKtAzJW5
OOd6fYNoQrFAx6bP2nR/vO6MUifVYpNpIgpm3ltZBSd0l/Rc5Yd+wgTVzmMen6Vjxla1PGdbvqAF
rjftdlZJoi/Tdvqvga4v5WHSGh56kMn/NtRC/ft/HZR48oN94B5AW1PaGA6apeJtbROscyxvEnqM
21PJn5blSqfI1V6j0Smv6FZlCjqwLnSLlYQkmdZCYk6Q8HXtZ2TjtJPJydWFa2QwPZl+UYB5Ss6m
PO8t8j/B8aUDVkeYiPWBJwO70x/B3PAylhsyGOTpmsMEb1IvolCw4gQQQg+L+5xKwV7DYlM8Qd7y
wwGxfnDGEe/BwbCDIWOA8Jg64sUtln05BW5AJwO735xNWNd3XK42hZTsGf1h8mQuVOZF3EGPXM4l
5NTv9srUTq7IkF1S87Mdf17EUj504faEqCuqogbg/udmooJJjP8FvdpKjnfNyug+XI4mvWoW2Hzf
w33sBDCPHy9Z12IC6ovh3rHrNhvB0CAk/cpnPsxkqua12pqhmcB748wHEoG9YpvSi0k82fWQ03mM
kOqBKLn5w/Yq+H3GEsBO8BFdIZk/OP7dUjCC+iAu/Cyc7MwC9Q/roTcdO2j2POogZRoFR6Bi3A2r
UZq1fLVIXgwvznTOBfCGs91uMp6KmU6HIHoG/QkDGfAv+nH2tKAT9iHn7kI4F6EvEj1am76uZk2R
lg5LDlqzBcPYqjMsDSWOPqRX62Jia2HQoGNZHB+JGndTX3OTYwLlT9PvyCiadWAO9pRgVWkReQm5
Yjq5ukfmNVqYYI+96mUCBKWNLIPGq4E6ezZvGO6qnonnzWP9hNZNKDM6eS5uz7Vd7WnPcI7QhiMd
17N+9aCqMa4fe870CYz4BsTlrzf5M/MxQmVb8CKRsOsD+m5NcboLHeNFS5sn//xirzx0On/fluDk
XQSBN64uNXQXuqRmVmRUmQlg9VNtN//RvwwL87xldYekUswjxQs8Op++lUNYsWbf9unYdVc8xGcC
n7Qdc5/FSBPYbaFGo/yr1tMt96VFlER58OKIVrmSvXkDxpl5Q+YqsOzZQ7qspDlNUN6Mwx0lSo9i
GJF8xzzL+YfUS4M9t4+BCjFaprd21McNibZve0exrIYMVHt1uFqLRfs40p/3cqoQLn4S9fteqnLC
0kMMqT6Hlo7LDIiL8JF1KPX+ZuEQfqwGM+b6GBd1WS3coTZ2k3JBKfcwxwDcOcfOYMDX4HfzwDCK
iZIqZ8/iwY3L7Ne9gmdlSF9sdLjrZ50HQ5G4PvnrC05S8WFJRL7q7u6y5STo+uFt/bT8Yb1IHOQC
YJKvAwBTH3SsaU8jofwDRrx8DXUngvlddixyC5Uc0oG50mQpoMveYRUapkfxXLZYnoEfk1TD3wj7
BFALHNG9Hexiz6EwJsLr84dql9FS39cczyBiLEt+z9psabJi71HDe/zGMAceTO6HThURoG4q6pPN
RaiyagkE2vfCRjGlb8gPCZuphkcaKV8kBxL+F/fvRODAQvljneinIjJBit0qPGfqJbULvLjZ+Fsh
ek4zlIOGigL7wpL63Pzxc2TRIYbo1oalSbCR0Wc9efGRByyBe3yCL+EZJX1Uuq0F9wHfJy2wndaL
6Eik4CG5q1SVxwivfKHC96hiX6w5c4x1lX39Hqfv9LLdv5gqOjozaGzbJF2ER1ByrE4T2o2TpPnS
R1rD3SbcZA0tC22wUYrBLYdfcPrTPDRKdPYmzx1NXEeLapN+4fviWarBtNNmZrq+U4Efax57oN2N
XVB/QxgXUC+xTH+qXY1GSo9trkmtLE7WBXStaP5Amc9C6bMRgn2YNqI8NLxyTS3ediwGrEbUE7Ua
qu0uHPOreluZ0yKUla7AkPxpI0c1b0rIi5GMp/SrCt4CdGVHgtiw6UPRLopcaKGUYzCeWpEAWrw+
vGq4INy3TclkQvpRXHAPzOxy3DmIT0D+GN+YISjIPe9c+iFocxDDhv7PlQBUUd/r/B//OQ4jDKqF
R9eVWIHiuzFr4yia1+CIIhopQ5S0lqhRRJ8NhSYKs1SwxWX6SRbGmAyklXv0rBdgswpvptTeoeae
vWPqrdQCULLM7PfRIfT0b+WCxf5SL/M5IwUx+pzlgol65g1LU7jVn98E0VbfZ3UiKiJgIjNEpIvP
38FIbADB5RfdPVVF7jQHPcJMkSleterkXBBPHbjjyjM+ICa3SL+RWz+TlI43pZCTmFR/uz/hop2Z
Q2jF/MVieY31Khv3+rXblwxiL8gB1qQF9C7ywIQ8Ltoy6/pjsGqLa1AZqWn3PRAHCXzEappoWtOR
bDayK4TWIxPBn9mCLkvONksqpIwceQd7DI5sK6AefvRg4Pq6pOqzYEkACJAl9r6mO+VWR5Y/TEC4
dyVuWVMHQEvB+GKZhUMnkU3K9euhMsVWTkklPbBzKFI0ifcAgnMnUseuw8TtLdsBcY8rwv4yEx0y
9tWFXuxKqSfho4nlE2KxZ/2XbEY2WSem5Y/wl92FG616uztFeHdShQmAg4WoHAcVQfkfszF/YSjJ
ccemNgzy5Hw8hoeWoot2V2GJ89Vv2aS7rgLjQnPf3QUZNGG+rcyNPmaNyUydm1mdJoFGO5A8Bijj
yZ3HzreXdD1Ad/1m9paPbFtnB+HWzNoJGp2MhmYIUv2+tQE14QYjHGQ1uerYC/YW8GluCzLSj+4s
W81OIwSnYBfaMb1yoBdXCSpURKeNCxZT4FwOIMZ7Vw4t9FY1/seayxHpSCIyqJrUK6WRCRc9Vwvf
00pqa0Pljkj9v184iaQGYUUrcNf4UOadxXyAxZb8t3TArqMIAJ6A78a5foeM0+EocJizMmgn3D68
HYKFBgiKqTmYnC6Aj3xjj9EZtQxaXUZZ4DyT9bSq8BKdIfi5PRm6OCla1z3fIB0FDeQRs5YsM212
MWGV80fiVYaBVCXxtKgG9P0CVE0MTwcq6xCo8jIuiR7CI7vHa/dWR1eDj9k1oBQ5XObNr4k4F4dr
tWVbYArbX4slQ/dFjlp2CawIZEaW9psSxGF3vfq4lJI7iNINAGJoyeUfoWGwvrwffQaCel2n96bA
27Vi7aS+G23gA/jGs1ZnbhKBtz3MWaCW5ztdXVRg+xFMzLUpQx5m/ULgBfSUZvGhEPNZyLVt0oxz
wXj6gVE7ybx9hUURXojHTcXosPiqBzYhGMc2o8JCT4gGF+t3E2q8YOMYbqWG6x/FW7/+/zA948rX
+nc9ED/DdSPavOXV3mT2WI85BIPXFnJ26a3TBF6oOu0+fa8R2g3njkEuZGl+b/WyAYkXU3KCpzA+
7kqqdAJT4+F72X8wcvohUSUk1ZpqFT1pCDAoLDmpTebwvBqn1v2UU3xKl75neTUhR8XiC+Vrg2af
tkE=
`pragma protect end_protected
