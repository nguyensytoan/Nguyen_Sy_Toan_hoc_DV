module  ram_over
(
		input [17:0] read_address,
		output logic [11:0] output_color
);

// mem has width of 4 bits and a total of 400 addresses
logic [3:0] mem [0:89960];

logic [11:0] pal [4:0];
assign pal[0] = 12'h000;
assign pal[1] = 12'hBCD;
assign pal[2] = 12'h03B;
assign pal[3] = 12'h888;
assign pal[4] = 12'h555;

assign output_color = pal[mem[read_address]];

initial
begin
	 $readmemh("C:/ece385/final_project/ECE385-HelperTools-master/PNG To Hex/On-Chip Memory/sprite_bytes/over.txt", mem);
end

endmodule