// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:32:03 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kMyMXa1bz9J8SLBd2dY0UQgj/gaf5JD7D4BeqICFslOU3MhOtSCQpfNPZ3woPpc4
WqnEGfOJdDoIOLu+rB290yij8YJ9PvqWWnN3p5G/3aRnVVVXiW/MM6QCS9n69+2X
kBuNtSBVLs/tes0bJ0dioFnlCoG+MN/1tfnNpYoffdE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17456)
JEBzB4QE9CIfuHyywqWumdJGjDIPpGMMTY5mwfpqbmSf9Y5TYiCsaLgd2dprZYSQ
oz2nksU1Sg4DGsuZh8EtakEw39M1ZytquzDmcr5USPEoXZvPvRDPuzWDLeLmYUVo
/YXQaRTQccXhc2mI4MTLT2Echs/N+gAQVMXpCi2fLvyThB6OS2RpH+H8pFP/a7vK
Dmw6IMmbHrkzrR9B8PSaTGe4PfwwSEETfIlpXnMPhKsqUSCWpjSjPtMDIsK7czfb
hxK+V9HuGr8eBllOWr5XizptJ2dqFYfbr8SdOUpxWwhDhFe/8CDPqxGzA/zTjn37
UXLz8zyweW+vV2MJis9n6HT+tm7gt+/r5zCHs9Dmp5GkZs/VScCzEq6O4Ur49KJ9
97gMPOT2224Vp2FoCoq31xvGKSFLfBP3RGg5TAK/N0Tr52EswKYYmIdv+32aTsog
oCuMFH12squan0WQmifnudalinrJLb32g8EZT/MZEYmNrsG8ssnTvnCfOoLQeaUX
NduXtefD8YvlGfqV5A+iFLEFvlwy9jqRV85mxuITnkigWNPJbWR19Jev7hswR42T
Qtg86Ffest/Rh+iRPdr9B157OzCqWLPdCf1Ulb3CWNfYWWzjQCMNig0GyQqtgyi/
57aT1KHp6PB7i32+q9p+fInCYRUoVuCJUSzeVOre6ouOo6+54LW9Szw91NAFVoqv
CNyDIOAIPRT5wYjM8iHSRh4Cx+7Jgq+J8JblqIoKqCsgljjztN/u8NZNY5hA89OM
5dHMGMJtCx37qGsaLhCth82w0X8NZZw20v/n9W1Zy6iN7TSoiSgP5a1h22xvh3Rs
t4DDLs5fDonele5IjqfCQ6MBSd1b3Levhm9qjI2ouWgYnh4t0muso6yccvDkzM0y
0ufiHpx/dL8jaGU1vYbKk3G3llbn5Gx6LOnlLJEsWnuW0PzTHi5cRPQ4OcLpYtOZ
r2BSTYCeQeDYGgGRbXN2MQKq0P/LKQD4jTV4AZeQO9dBa6PpDKRhuCBp1kbN4U+c
DRLzFGxP8HfCQE+0kngwsyaqHSUFSEuJIxshyUbNmr0loNfKIbsIZFRbNArVf7bt
MsxPBF0hH8y9h4CB4sQC0L66J3xIM606NxpIuTn0UpCOmhjF4kEJjyA5n6y1/0fW
XL7EoXBT6kErWs9v5CGhM4kzYYVYmkl8MfhmKHmDjfEgFp4R+mknqRavPgb1QIYr
q+sgWGQlHR967xIJTNnE731Md9wsIwqzfEtJ1lOtDXVqb3mf94Sj88hKpc9dp1Z+
WQE+ILyeH8gjnHnY1/kg86HA4lF/ZtWVYizYg1oVvsiedFcCAcK14OSN0WH8V8DC
6dP5Avn8Nfjqyzlbq3ok+WIJH7NXZAsXWaGC6YLQAEjJr7TyEtb9lar4qWWoXQ7m
ibUS5grofdRZRdqFVxiX3SOnfOMb3OXtSElOHRzD+aOxmvodKYSZlOeo1VJJ93DP
+km3pGXlPLkO2W5f43fFYY/3dyNr0tyF5nMQAdENY82J/gc5aiSKihF7+7GqBcSo
XGVJ079JPWKPYlni2csPz2FPXqkzVy6aKEoNl+u8yBC9J9PITPQgBnhP5Dld5h7K
d7EyiQEMeFYTgXRHIdhoCASMiYU0D1DmYnf2gjnFvwKO92zftIb7+4plwAwbvPbM
I1vFFHBmdnxGYTsW8nxNrkl6ASlzTa0iJwtdwNdUUYDdw3aXjky+KFu8c4gPjDii
LUdSXyaIYAhk/lmj+HupUtTDZHYEHq+odKsjuWI8uub1GpcVtAagTY4nosJX1bEZ
MgheNmKCHuz9tAqVBtWfGLvQ80LYPLCXV5lkXbsWr12CV/gytz/VZetcQFEfPUN+
wAZEwdCbjJXflfWt0FYDfrJxh3x+Z0W9q4Hc+SzCzn13hktaLI+60zUdieRx/8eR
f9iij3+QDgVZYaV7tpKuKVDShny4ZL6fBne7zHAq8qfXaojxNjvMueHUKkwpbsd+
RNjG4Xn6TkuBvFENxMUpptbPRfbUrhhupu9O2ajIwf9vetjt3jgzOrGqR3xwjZWZ
U8Pnsqdwb0BeAM1pZTRhRVGJmavAEPYGUnQxkuCDjy+l1NmQg7maQE1GWum7HsTR
umIdMCfMngeQ55AddjhhFih0JqnRE2/OYMVhsLE0Mw6ftaWIr6WAKnunIg5OkpGu
8LZizeQaTYy0+Ad3dwCn8fwBXfpKmB7K3k4aXfvfAOw6ldHC0hrcnAQODYMzXurt
boRyaoL1ECbk8moUfzg/bYSB5rrodCsay3X/w2RMG/EG7nLD/cY/TUhLjSQZ700+
bKKQNBSKdrL2afk4L2aT1Ok/4NAZuUij295a5Y8QsqvbUcUIfqvqR4e9/KBc0kk5
C9NZuZhawemDyVoZYZx9M9jTjkEa1kz+QJckRDSVT4utwo+aW8zooewj52wCx9+/
NS9azH5DuM/WrXiKn8ivFmeAU7VEfCeIqRxqZvbbq5LGgIMzRRuHq1DRq4TAuRdJ
BB7bWuU+30IHwNzdKSw422B6sXZQQkOkdGDLc5DIrCgbf1eX+ZBrA8Q9EKAl6Yjo
Km65dAg1Yy4DKS5P3qEWE1qxJUEHNe59MrGpKo7OnesKOTM6Z4c/lHKCWekeCH8P
jSKv65YKZRVQhq2IB7r4/lGOr6tD2yS+CM91Q4uBPUHKTfHHL594gr3CuwzNmMbo
8a5zGCZFwaohGbO5p1eTAAfB1WntSB0LV7kxKxhJW+N3jeQK/QPSdiPMI0gJB5+b
dDqPiog7aQkurNw4sq3ZepYtk7lrbqPDaL/Jgq3D9vAYmjT78AP7Tni4LdivBTfv
nnxShiYzfnnwq/EZJcCWubmccawjnwkyC5/b399MD3WcumJ/jRfXMAEhgboTWvFZ
3WTprXwucfI9D+itXRUWwkky2JIhRsxVHMKVKU9l8/PDRkBMQx500J0RdSU9YkHz
R6O2IlDPsJl3mQU4j/AnU3aZHfn4hr1A7Bh/laDGlqFHcz9P6dFdvf0zQFMfY2Mz
+9WhyvkeC7vuwoHs92oaMsIwt+ngh4C9nCPe5CYNOg8Z/SMAbKLWanAG4KQeb/Lc
qvi5j0JmPQZmD4RcPzTSA8AFi2i6rH9pvan+41dQF3TTnj1UdugBEGJjd9gf6Sy0
j0EQy/gndiCSFVX9ra2mpoGk6ETRwYLSjjxiMVu4MOAAsRutW0SdHrBck3UjAc1A
LS5X01LiD1PxeeyLcrSDZ6rGQu0gIit0H9uNzBmS1xYsGLLAw3RovXYevDnwviK/
6EAzXAZUYXneFYjZO/AFZ8lUJoEjKfj4yJsPOtwX+ptXyw2SNG+YQjg1h5VOX+bZ
2YWcoKw28M7C37ITN8g4oV1q6R4mAqAIVoL1mJ4h0JF6Z+robZzlixl32huEK5+R
O44y0uJ2YPcCM+pRkJ1vdtauKD/v6lfcE0ASYIWkpa2yVWN1nbIj8pFWHb5ckQ1x
pVsDZbbayTA8lfwR8u4l2LxGPJMwrxhVE3KAt1ShNDTDfqkucH3ptOll0UvLN7n8
j09+0qC+fshCtJG3ZtZGD7h6GkqQEtiZ2v56GWn8PZVfKHftnlLZvqmeI+OpjxgY
8h3ThrkqjXgpUiNN8Xw1f24kmdPR6ovGsOojDT1gR5sAj0NIfXxw8dexjCOVDKRK
hxcQl9hL0KrU4a/erGD+eWexJlIse5VSP7QIShv7rQHITK4eSsqjNRj0NTg4b6T9
oZP/WeP3bi2hD/z0UQxlY47+o1RYcKOf86ln/9Ev9FN4rQ5GbwWNvUJI1SJECdAp
vPGBlFx4Sb7yQg5DLZgIfVO2DbzV9Y1tenGn+zXV5QdtFZkHdY0n10okN2KJvlrp
zs1QdoLUfPt9ld8DAeZD3Gybl/PrV3chWOPL7+fC5jXbmi1sSZc26X9M6RPF4ELs
FFWZhfQqGGQ42VMMMUU1uL7yVHbutq/csZuEUcZDY2wuAp1KizGtK4YzdAoXOj0g
ZAwOWUiRSt1w/TS3L+k8Lluw0UOa2rwrXGNvzC/UPOkxPl24cWhUURW07BacFIZC
Ix1+EoiDgnboZNIPrBLYBLFVJkJDj2zGM+33p71ZBGyB9Tu4OaJqMCSH3dgx9sRK
ac8rAxzd2KlaT9cTtvaDCt4SfKMEWKxJMSO3I1ciGIn30kYO9RAjHaEWsEOw7nkT
Pa/g/DM+0yk/66zCOy1L38iOEhJgr8TEIvwq8bHswPjub0YNFsQ0JxW7zGRjINBN
1UDKoT1kAqy7szLIWCc6ga/SU4OCqcde0Xf1sjY3ztO0H2R8K6b1KnWcp8fFL/hp
h+hYVWL7mZLz1ZPlnM0m0d1qk/qJNA2Cmn9nXY/HOixaSbKI7jI6pnIBJBGN3r3K
Jig/j/ieunbb2vQ7ZcarrK9ClJFTdGEKb1D9Rh/R4AljK7mRRaIJ0phU1C6Ez/4C
P6vnSyBbIqMhkoMEfEAjJUxqor0gh9kZ3kDpXwrdbVRIzK0s1JKssFvXVUd7Vc/p
J0MQiobNWzfHU1IlWUcqoLmqcfMvAzbr6j9rvqDvy20zOGs6fplorsxBY5DzJKVd
jvR97BT8r4c3TDbVvJnd2siMNxQZu5OUXSgeNNUcHyyGqsluY74DfX5iIuBdxozf
fq2EWlB1OVfY7YO4BfLKZRiAC1fviQ+lNtbr6m7Set1zVB+GzAjtRiKQhr0+GOkP
/4z0V+NO+XaaTxA3rnCsg0W97X9NgNt8pt+Hg6lpY3LWVCcap079N3q/gkbQWgzj
eiHDOumQL2Oneq+WvJEiTakuTNLqJpGHOfvOs4LlUA7pcXLf1rX24dWK/FstXlRZ
1Xngs3YJvsddJNUvktwblw4y2Q6jioT1Pej7iZ+bETz/zecL1GDK0uCwrKK+RL5q
d3q5towquEVsFgtEJofshYh6BeCC5+tgyiAQ2uME75kvpLFYejvgU9azY042zVAX
R6peB37lg1nQbjEJdOcI87cCewJWG/5h0SpzgsptZDxhlxGxl0fL6wPKgHrxT90V
rdrab2oyz/uZXEr3RIGJVuZ/j5Fzx4eWvME4PdvMcdtPG3d4zeM1YuXAlFxaqeNQ
BhiasSkiuuezYgNY4GFJADWriOr5JEvqnFUkCm4lnRt3evrtiwEDUfTFqenpVVxp
7tnna3JoREtGrl0JEbQn5T7SGUSjbyCI+HtwNPzyC2/bmELmXERIudP47gPaV0Vx
dg5X7G8K+gAK1C8O7sfIRKG5lXnbQMZrNvMf/Ee6KsYMJom1mNGP4gxZIJ/8T777
LJBuuEJ8XM1Ka+tAzvqdArRkTfcUOJVeguMUePs3h3rXpGcV4BqA8cuiqnlceMe7
Ukrxfr55T8FTZKKT4rW0wVrEidUJ42ra4jos4B2zc6WOzTPhQ6EZKVtCDdRjYQCZ
j+Ui9tfJwLMgMeITY64YujNvTBIpOluI0ZaDBKp/h1epOHRBFu77zDufQgSdoiNr
7XJLlHau/GdKNOEUmrGmSnOrDoJW0czv7r45qRGE2unmcBDZTC8SQRPbY0tJMMIJ
dV98e29wLzPRw8deOBXyLldg5xLf2411bEBlkoRUPytdoGilXt1CPFd4ARtwL+kA
FzAAlCqKKhxm2scahc+Qzp16akrhdLJldCXE9YBkSUnPGabBdjEG34Aud1all7Cd
xLuih+vRSPy+X4mHXwhIAsIvRMmngnmJeioGhVIwUQXoDDxUuyLVACMiobxWf84U
zEQG2BfMHZu0FFWG01Y5ITs9O2MEwklXkMX8DMfwH8CPwx+XEny3azbvsZHKAavY
4X3SnRB7G/AFYuAO/DrobqeCGRhUjUvNgntssnJtqwxxxtUNxDiC8SVoRIcYwmRd
h9yiYe8Y3azh5DPNcePTlrbOrPWx8o1OH8s665k6Qfy50Nc9N7xrzG2DLDWDIMFS
vJ9LP4RQ8LxMLBnNXE7nh1j3thgxVBCW3kGQqq4coi5bfUF3vjIhUWvr4HlnerdB
apl1sXAbT2/p3tpo3QKV4Qhvq1PR3VVCsjnM4SVhiZxiWoq3gm7AvbCFil6d95/G
FrSqTL8n4/wRFXWYYeOFpLvzlYJuWAWIVRvxGzJ/SSr6vWulBCv97gqHnWM0iM6K
ITI2nTO6bjhjN3vucGN61u1fnBuhqnKNNXyNkquv3V3GhgTop3o/47ODyLA18960
+u4tSwAFPdtAhxJOm8lSevZM+UzHMDuD134BUXpvo+ORZiZypxE2AlCQj+pLbNCw
Jkhr7eN1Sr40BAElKPHWLSlkcDcTope+WaLsX+Mi7Es7u1g1BjA1hmperfGJAylo
vFLrHvE+EOH9Q1RFURTbF7CgKSsLM/Qz4QaAL9STyMAG7Ie0aXWu6knsT5X7OXiH
ezoRO4wtB8naDJiTZB1jUVkWVj1aZD5QoSGzkgePH2KCfcZfBHnXAldSntg6BMKw
SGF/77osOs1KN4TIicD/W4PxPCEJ50dW7BX6hM1bCsa92atf8lE/5iAiTOVpqJA6
fhJDosJa0wLwgUTErHXIeudvPYYHKp2dTBZ3xMGi8+JWpKJ7ZXJCAJZzpZEbJBcL
5cQ1M9tBuqLdx8ODcCNdUd5znJg5VzNyEi+sX8PB57SMTjcDW3MHfeGYqkdrEab+
TFPH0HHhKVdt0csn/RHogxeGBHLpaXhumRjWxTlWXjFpSzub+AOvvtTGlzjJbMgT
RsWzrgHAWEzRObFhPuUeDUXf12Q3YXZyQIl9wMyU9mDmxcqt54bf0JVEJrGMYLjA
nyvYDlLI02YJMeviwNZ+1YA9m7yJFgDDfooynz9e6jRCGfgJ3GmfCBu1/tQWEcTN
dxBx5OZA11X+te4qjlhpo8q93dUCY4IG3BEwzSmI/NL7TuKMygEOQ+nXuwWhXbIu
BM5IuZu4j72eCnx+oFecOCtbfA6e0jBDX3xO1rlEzmGWCmd4tfuQTCTQ2dIjG4M/
ohWQ1mVJOI37d8MXurZtjM51w7cMfeoCEXTmcTb9B4nASy/Gm1cLyHXZHvXDOneJ
bjW+Wb5FkinLBZ3uO05R6sS1i4OnCSeGjn5O7XwpuVCHVLMA1MibFgi5r5sEVVNc
Z7G9rxJvgWWge4dyQU0qR5xJRN15YwZzcWBUrqF3fiUKhbDWIJHNEwZl9ZWdGsaz
3BoGqwSUbtMfJru9kVxIqRrMFSuRy37OXG6nd9N2OYF1Ctu9NERSgKubFfYLCWFg
+QdtWk62v8gGKjY0pG7rTbtyVzW8M9GuloWYPyS+qfWCQ1lcKY8GvXuzeK1ccF0a
k20w0zmRllmBEADCP2YISGbhCwQE+03BMUtP3C4S85/0JdHCJx0Wrz11ThvbbGAd
4ptoG+tjVnW5I3cHyKsVCIt6fom547d8aL6D8gR86WUVPbBkAvGZ0/AUEXU3pdMA
uZCVzN2iJZbKxzwoC9UIg7SO7AN/TG8OqYJRrQIrIhrD9jKV2qNYWJPFkNOMPn3r
wo3ZAveojw90hxJjNcA/HvS8yGr49Fh+Mb6pPRYtUTxqa0awpqkCmR1aD6SVPw4+
jqLd+e/RZN9IyAgmLRXIdtzXj6sLEDymZcMUkKnj0YL2IEt1FVjGgg/36+5ODAD1
w1ZJb4/7XVJD/SfMtth5UQCcSPeVCFsnN5DDWwpg1B3clVxDJIPUklMUX/zXFbKQ
nr2jJGEwT6JwKDJQUfC0Otax0StfdiV45xTScNJV6+fmEPkOZlcqAbLaz13JEBSf
n1F/fnkUpex2xu6nYC9tLTj1lVAP/wsK71Fu1os5vruA7k2uygJ0kyxEEOg/BW3z
EnsU64L+ENwQa5Ewyr3fhg1z6qMucZeBJtjdFZVWqHmmDUesL0RsolJX989sYB08
VXf6EPrZ3tYDX8ScSKf+xCCIgx4s0Php2VJ2C9Sqa0RHtovQJoCqGzAFNiTZoYZP
CbGGI22tBZ12yful/qWMoMT2QgJTglNeQxKXwYENMXXHIt9uKGo2rkcCaWFbtm7K
wc5vgFkS9zjAu0oahJITzeivYD5E40gDlsw/xemyJOiScaThOn7K7RUqinq2xeMV
ENrqJuxSUQDZXmDNycVzEQn86KgkyA+/1ag2Ipxm+EtpzxSkOQqeTaWLHju7K+cx
YCLY6j6G2TQUPoLBJbssWYiWm14sH5TBd8e9Y5AYe2w9AZz5PEKsatS0LEkqRCXE
tWmO7C3FyKY6q4Zn3J/gkyCD48JVILFx8c5NcgzRFSFyJY7s1BS2GMYb9R1DE0dV
rZnTXUMupmEM5zU6nhTTem/ocUzAGHqPcSvzFRxrao+47BW95H7ars3Rvkr+f7c0
59y9D68j1zi888UbLetxsiKm0Dngjgs0J0pPsJbwrw4xj3xY0MsYM1/t2nffuh1g
ZuzgAjxY9OjgGA9ueKwybmSWUUx+DyAFdWR20aBvs9NWyVEiCqba3ou6qsGpnW+I
YmCqEJtLQV24pO8pZwu95vTWw5mvuGEreNbSPUGl+/v/0OHuXqPTMhorarRie2lO
fGKO4MdMk3pY1Yo3Y8draCza7WByDvxm1axsERes5pR3i+0+dkDtlRTHv3qNWojQ
wiCOqKAkuv0zoFftpLkrJv5nqSNuXcK9N2RS37D2tJVNkSOuRS6gI9uHsgSKXk3t
6/7HHUY6Or8QSmzVxbRu6wexDcXp+mDTFrGAE9Z8A4SyBXDtwIuDiTatSyHeNnR5
565OfLKH9W6eEERBZ17gka2KrAgrhZh7ZVA02AG3nZaNCpSvcryYJRwhsS6VO5S+
IvOqYBMCmaDVpnoGxjY48xD+r/tEMr78aYW4r1eyAxqgsdocqlfhF7ESOr6gTGEx
V99MbeF9pEBPfJv4E7OLoJ0j2dUsatqjtm2QiwTcJKRMOeosDIIwbrB7J3Io9UsG
he+CNJrTVNDCMJc4WpGy1Jdz9PE36+Ptil2IL4xchUGyA6xUXh71LX4uwbMVXti2
NJ9LRVxUUPW/OKKUWQLeXYJEx6GqjPIXL3vCFaaNpx8iBZpYWhvJPyVh9OfH/Zuf
uSzx/WnO6U78P3YaxZ6DuhOG3Wh2UK8fS5FmLpfeUGMNfyG2uMI+cpcj7sLQ/+p/
vvhzeHkSJ1TUDoWTXkOE7xQ/1x59rhnRhxdGFskdH+c30pYWQrgn4x3BiAslOZ+q
IbnapfFLna6zeVobFhrXMVml/Bi05jjQ6bkqNUntidA7YBl9wBUOifxBzGFXNzUj
YlON3RZ4RCx7uMJQXhiHmdiAQ1B6tP6I6k3OvG8bjqs9oCMjzsy3vDEs2tZNGlNM
cbJdHeywdKhyTpMiMNVUGSVr6+pIuRc1dtbT1vEiwO3Hhy8Fnhrm0abMYf4tHpd5
/f/4y02gkdYNIkJdStVcOKzO93KyewRoBI2MSB6yJW++jwhQeySworUmUBpt3O+T
YdeqErERJNhNac+EcyB5tciUrtLulqDkynhpoh0Kh5PDKi83fU/74QvYTVxmCCBS
/n9K0XUwyhvQCe3jkbWWuh8WztyQ5m4DnV6zfc207w5KMZeiTsh3zhMerXpDwxNO
rMpnEhxPCTXm6QHuM1ghtoeWevaIMy6f7ERB3BYX8bJOoyxM0ySU7xr/1Xz+GFfA
Flb+2BVAFfvkZMpOo2xmh4STLreVypTSGjASMyHVHwYM06QTocIOPiW0la7ZQHsS
Cqki7+h0RLsFCxdY2GpsSmXArtxX+63LHRq/Wbru7bb69prXRFbyLXO7S3oB2hVI
AS1D7IuyNHuKQCjSrMJ6Ar1jetEFdV3LnTTJclDF0Xhs5WPS47HLfvKBv+zySlhB
E7q2JRiNjMPdi7FyCdvqdKAyeLczclCk5tkdXdip2qSpflx9GzgxvgnjyswvWRPR
BI7YBkmWj+92RRM1mH58iknslTQRE00p5vWJzqVY4/OroNonRdQhkdUksT/61yge
ohbY+HyGo6kG5IvWZmLPn5MJx6NxiEuaZxvdU/ASrv0xdc8Pfm9/FHh5DINnOjZp
kpS1wraoMpaiFvTkFYWRsk9N3fjXoNrypedYCe4Mv8YMlfOrLzMoTtuVcMrD7Suf
figsdPc1nfxCRLqnvCnaWDmcF4ZfAb1Qr0HrGcQdY0MzlDSiljdFc3bpNMy6ItKY
rinmJIongJnqX+Zhp9JNvOxtOTw9E6YZTWHT18aNuARfOxw4JaQxzGtfN7oCcfTO
SxcJiQDKk08atRVpIlwikQNDdv2riiGEeJGpYGF22QiHoECHLpBtWpFLUj0HnHtc
XcyDwW3ZHdh9Lgj+AKbAXpX8s+HWq4JklxU+uLJ6j6MA2ssgK/NyvkQfqjMS1+Oz
0mziXYDG//TFmV/Yl7KrcQ5K721S2+98B4JVfdzYP4D31gCdwzGM4O1iwjPTSPVz
taVT2g/SQzpE4Lm/ehdmFtcUBdPEyYKPpAa7PXGmDnG9MEaKfxky3oCZE/4GymGh
dTb0EOs6+IGlWuqAcMuEvpdnMjoR1iR/0PTS5My6nsNI1FFGntjH//fr35ONPPZt
MuaK5M/FfDM0YhCwzwJtDEDbqC10hYEKxWKwpSOXjRE0+jeqYvUkdw1E1jmvEFvn
JDe0MPhBNp9d+BE9vZoKIrNPqvEdQaIUAajdHf3dbXvlcXvbu6E0qJlTXb56r3hr
J3aIyckVVsr+tg4oe6qQOnITHpO0FstmkleZpz2trmMJJT6FiUFefw8DQWRbqXqa
gIZhBe9OUoqo5P8TOchAWHF+pqerbDVqvMEnI2a/5SsIIc8hiJBFoD6Zzc7FSmNg
Qwgl2tREegBHbEthXMmoLGZEVDNPD1g3/Z4xp/FK3m3YN1fNsu2iUAKP9Q2zRDyk
JlLbT3tSv+g65WnHcTDIwPsNmk0Ag9yUVvCTGT7R8J7Xz7SKUdkUqiMyju4U10XQ
7j/tw34m59OFVNgvNKsDcvEHjF3Bmt9Ta+sxdXsumo+QyyoJBUCVycpd9IlZnrZJ
bfrDOQB0BQ5gPYLMWwQ3H5e+iQ/FdBIEYWTgzVAWNvzEs/sehOGy/ieV2Ptz+OyK
iL7Z+qFglyUpllLQqsS+kzCklbHRgxvq1TCXMGXG35NV+hPV1fy5gZBRmK/tn5as
RSskDr/UcFyi/XdEnsrOhEWwA+ecCpF+QWsHhIVg8fG3BqemQ6PPksmcVW+2XSWu
+am1w7HK2V3lu3TGlVm/HLSDU7MxULV3y99NgiuMCHZ4VZxIkFZYZmdHAdBtE93L
pEiml05llqd7+xJEf2ehrG+sov5ChYIxyEsHVdN27voKIcvzTQD2Y0qWpnwO5Wn5
h1YeJjb3yGZhUQ+ZzcCsCYGaaK/9A+XkH31rLzzCy2ziTRFIUR6Thz8nP7lN1JxJ
hX1NgUZmJEdIlG4R9H/adG2QqXVd09xuM70OBmQb5sFMDKhMcgC0UvmWNVnqFTB5
K0qH37JnJoQXRFRvMCRUQ46wBPPUapIA4Njfp2q2XdEI+hGCltcAuSLrnffgGvmt
Z+O6KK+siN10447Etrf7DkZayKwUfFTrw11sbtiPY3463M1RTXk6IQQsvuoADutp
xVFF2k1jE7wh9IS2tBiHhG8ZNOgVsJQCFqhEHPp092m/DIsUvqN4ThI3KQhJnCCP
/4KgpcHou5a5ybndx3Z+UJeI2s1F1XgFT/8GlDAcod4gPMf+Z568dAv6ac0HkQ19
JkH5Hcot03ab52X7qw3cMFUicJqIF7lt363spGA5amP91StGZQp4441Bq4Se/JUT
JnuT3uY4wRxD19q335ol5q3EcIAc7JXJHBUA5P9gcGZ1OIQeHLqiAZXHbJn2QUtG
kFXx/UCcl/657cS9z91WPlEk2sykaWUuBUVj6vnG3vYfRrE+ZkSbGIWrJtzgkN2F
TGTfvXrHD8CqN/TuO1di+VjfQM+qEazoxrwa4WCn19X5/HjHsQ6iiFu7VCN0jgit
kWABerkDNfGPKSR2nfXYA3g9/BwLd+6QFgxt2wdgUwF1aKQT9A+0LHlseDZn9QXz
IZZ1+78OOIp1C9Ppf7IdXPWtDfptrq/94Ey0XIb4rsFku14ll4f+WZgHePt+uLo+
ZpNiNSMS5LCj7njSGTMfHZ/J8y7O4GovC9ztUBVeLCQk9/9/EFCn8kIg8h+pYUca
l9upApT88m8KspNoxyb5uNGILNzjgIrWoBqLcMxLp6Q+7U1Z1Xf9lC7cNYszUS4e
Sl1UGnu3iI6ePT4+tF3YEN9/n2BI18mGcwsjPTzcriY06hn93ooj1bb/D4+OLq5v
HZ6/sVZPtHocwHO4jsWMsm0iqipjinrK90H4AooqtxyuTUiOo4XCgKBvFIvQ/mES
2FqBlLDpm9kjWKGGlvEEOHsCRITB+nCVz5eFK5rWpwAhVKKN3WGis4dTUQY8Kmf8
6oqW6TooxiGQXms9jlnw7XvWu12m/a5zhvVUIgPfrj6AqGv+sJIQ67BWMZAh7/JL
0tnG5kk8gBJFsqScaxTQPX6rHq7qEKxmsBX8qAeRjhJK7nAGWhaZvQM2ijAyba8x
VzJ0x48GQUsblPtzU6jE++WPA2dNxqPxHKtjFSO1bC3IbmZtgg1TNPeyF9k5zdzS
Zlg9PWxKE6qRUo09EcLB5qIe715rUJ97soTNlT8uQDoHRtxycfohgO5kyxi6n5gS
s+7olEgsrNGdtJJ6EjOb7lWLH4lQ27OLMj8Lxtwdgk1kQPFmeZ/FN1CZvgP1/5Ef
OuDoaFkwj5VE9VMHtVIali+nFaa6pwaEuJRNMuwQ3Gv7LO8CB1ISGQz2qiJZVtVt
/3fRTT7KOdhPsHPjD0xV0DNDA/5i3QviZby+4/Wl9E12Lwc7CSkikfJl1bA0J6/6
Hcq49H4eaVIeTW25DhamUIu2BCYgef1cOEwRWQ6rKT/h14Pkc5B7nJdaEsKL7X0T
vVlHOoFsa48jMeR43s4feGZqG1q4wV3U6mknwo0I2HtETBaf+VQthEkKM4vWi4qI
mInrjiiFQ+mdl4hOn6h2JrWOOI+gs/FkszJEhLM2XgF4/nL5wfwGTx5OHA5Sogwq
ziyBWYNbODTqce2nCXTQLK98UasIVH8Cg3Wu4K/m1DO2G+LLvxVfRG4BTIQW+qx9
cMqmzB/tpOQre5OqoIcCL532u2K/hpbdrJMaeUj6fRT168gOZs5f64QgyeqZkK3L
BZPHw1PeJElUoEBg/Uio6CGv/kp1AZUid/zCbJ4peQ+jlL1EgELUnfo5ep0CnbJ5
RQ6GxZZXGU0Gvycunzvfo96sz3oDM6NWUBeIjStyN/1GpmI0aO6RE5EZhjG9YoGU
Hfi8urcpY6UdOpR/8NB8nkKm/JREO49khDIyAXCLew/GZgqL9faR7RZ9RWqEzWuX
b1gK7BSQ/gxUtuIP0mazGscWaCMANBpfV9RMqtusK409GX3vv+cFAgvUu1nkEVVI
Fi/X1n5E8BiQ4eP5Ai17pd4lowq6uzfLKpsQeAZGApXB3JreHnIHzqAbRHPc2JgO
XyEL5Nj8HT5ch39XTVtzsv+R/RWd0tt+cX+6MfAJi8Ig4nDsK17wxHT8+OQJ06Wz
cqPeivumVxRI73lQ++jtFqUmcUPRNm2He1VWa1hQ1Z8zsh+UXVceEbqwwjoHvpk2
y9ymyUS4MjZ/pXqAN2ABcjWDUNE2z+Wlfpa2zmM9kU1y+7cuz1X9A0M9mM1nQqxw
02azWqYXmRpgpf2Cx/3X0/+wWihc8mB6T47hRy//UDlE3vecaGwRFIuF3n6w5eeE
nnuVYbu4nBCFp08OtxZMLYFnnQvSgdDfpKaR22F6TLjV5+eKLWbeimNQ/Uel6b+h
bYyAava35K9uto/pAKwTECPAvrFF7GGFlwmWu6U/cifeUNy4FCkyRMA5Cm0YlgNZ
fBQ00M1aLTuUhplKAWMvYLWl8TkQFqcMQ73YktIvWt35b30ngkWsSxxId2KS73GW
Zaeow3fCMZfVZTa3LzXr+keEIhe7EbHpmTqbNqM94+jVyWxF9As0HSFeB/IC6ARQ
F39b06jSh6Qm4CB3Xns9kQRVkBR36NRTK4+Hav7+OqO58XEUc97uJWbEwUxbWyTk
oFh02fkOpljJ3coBywEgtUmT2j3PzltSqamvyePVmPKh5PUUgXXeUD+7ong2mjN5
aLwwkYOIoeZdJr754DGia4pdcn+ooHXN/LITclWKSGN386Sc6sna0NIb4vnawJTD
jeZ2qsUF9urlSdERVj903IJ4mOizHrtnvXTAatNLObfH9ksFm81OS0MOOOUs+sfH
1SZJ4V6oMShmzLCvSwtYosYvRmk4bAlnoQfzTPUP6e0RduG+z1YZ/G37/LdEnHnf
I89CFbAnlgjWRW3O7xlSjazcp4KStTcrWOvAOBia6AW0+0s9KAvprQRsbEgszjIu
mCLpymCMjZrlrbsUPc5oM9Y1j2oiGLddW+8JqrVIKTypxN6c66XvVuBNEg+reNXF
eS0VGqJ+TqUF0sXDYuPR/DwFF/SqY7EzNzJkA1FcKapt9m8D2IuEXZN9NrQ45NTw
u8Mo6ky+ifyIUYqh7fxKYWeH8cJ9Jna+Qrto2XHa2DoYlFpLXBQtBzJAFuZyjq03
50/n4THMaHn42QHXtUK6IihaxsklKsbT8UxmFyQuDCdQQ8tzI279H5mdvn606DmI
JDGG4AfjvaQzmxhbTaA22nnVVxHjpBc8DHo1w+t8HUP30O7OXdvLRxhzIv5JxHxP
Wiw2wVRB+jmI806rd7BzKqkJp9/bmT9q7NSoDE/m5cGngOoOkvjMYV9juz3JqUjS
UHCHX06SqIgOsw1em1rVGoFRgM1VohMLanB6LszDtVXEwnpCJLFSOkvJNJJcMdjk
jbWvVXlq7c1w9LDpFaTvXrH3MOJN4+Q8OcxX1YLhbbIboLq7EbEpiHdr7GMLUP4g
Y4tQrILt5K+QcZGWia4OB2Rcy5BuCgmNmemCrKVGp/JTAg/zE7YEHi8OPXkdTeTT
A99DjwdIbuld5cCt93WiiCeg/51THmtT6W2qqbcYYwu2K8DCr/CnbQYzkWtg7hxH
QGoZiN6HS/B2FrOCBypgnilXHMs2WABnMifGz4qE4mWle73Vg+vEUZIFwRzqyJil
jnKo50x7b4KpigBJUyu2M4SqesmBZDTaRVt7OpuRVbAbUOEHTPnGN2olKCZH8zZl
LwCFaE/lNcrOnqwQT/l6uk8jmhcF2GAeXp/PZkRRFDuXwV/LlUeESHHQfmGLRT+X
Sc2rjkkjuR1SIih/QloD1IafibQcj4jBcGCsKl+XUnf8sBTFymVfvXqJzT7vXOi8
tGW55lwGA9QdkP0JHByzIZFRI4ZgMYuxYFsWotSm+ZCwAbGrkJMILo1tfe2XZDNF
5+oHlIjGFt9DKF3bnO3o5nwLWHzuMBPewYj6k30ZycCzxtO+vRM5rYxlsaSYz7wX
EqY/DbEohcWeGis7pJ2ra3ITcoE/0IwgRTp8dNS9irUIe3X1zG18z0LDB0VktBql
8lzq57YMKx0+JX649z981e6Ymbhw75g3u+/eGUIXvHjxXaLCHlYXA8t9dJVOrTVv
5DVXsap02+exdPHvhjeSu/OVvDZM3U0OycAveXpMHZ8HiqIPDDPYDpbsB4AJhErE
IENBjeqwRaSPMddJeR5dAkqH16V2Bk6G0qM7O068+bKBlHR17L7V8mdNxsvJGDDx
Kq/54ffUJVGs9BvPQ451YkIhePfUG2KUSQWw7KiLtZlH/Jr+keaH8SsZ/zxn7av3
iJFlBi2k1qQVbJVDMHPXirMiUYZeaSrlFkllxKKyX4T6Rn+ig7ZaIe+u8E7muSOa
1XGEaBdaIALR+4DcwPYp3tnA1eXsE3stxDsWfbRc49UmRfTJwhLWUnIBkkAxqxdl
6+OSeRsc3Hy0OnG4GI5ZUQH0ic3y1LbcCCxdaQD98DzpwbWi+Zc1x4z4DOTXOuFp
xc0ggw8KWcaybp7+O+6xzfTXZd1CePA6horUQnurg1cjEtES25YWG47KvY66X8GC
UmxKsyjb9eZ7kEZqyN8xezqr6TVLinf2xwyEVGbhoeBuVSK7oD/G2+qNuXkXhs0y
sFv38P7PZnnl987NLZ+TadS/f+XJEFGEkgVThZIJ/ErLQ7xFWmXx63VaPA5rDcta
EEWydQWEbgrj8bxeacErgelGWjwyCDKyUHWWjmuCy6l4JlLAgTHUl8PF6ox7kGuI
LF4K18J+8Ty62M/j/3GvC+c6mEcElppqjTbAeC/xqxWcO/+tdb1C+EtiF5Kfohm7
lt+CB31r5j5E50fo54mZ2GDaL2eBWK0DRzpSybKN2MYu/pKiQ2f8frxwSRTjfj+Z
HnHLzUfAxFwTUPk5kWMoXhB1vn67Vyt6B2lH+tuG7y3P45Nj9SLQTjFFBaIqO1eL
kqS29cIxwwuKesgM4UhyZF2nI6/xGv1HxRHJk09eG37F4HJ2MHtO81UVjQ0aEB/n
ZiDmu5wT6qOHT0TRedkYK+QR9htAQEvgcxESOjbHimcwQwc34JwX60ZYQOzXVSwv
cfsBg7EWY4wltMalWmo60IRl7BKow9YBPcNcX+kU9aecOm1wAONHDk5yaHN5SlEN
6Wi1SIIJyIouH3pYsRIfCLDwvstWB2pBYzfzKTx5ruyunPPXACr8XGTKy98H4t/f
hkhceL3MQBYHHzOCpF2B68M9CVHJrt46Q3jv40KyjdyCGC/LlE9VUvvoBUFs94kJ
kG5gaJzUEa553WQt/FdCDMrVhJAL0SYpZPD3hDbZfymnnoVOekiXBZNBime0SiKo
k/G2aojkSNcz9ByPSpnRi0OsIiLvMzV1jI5A4SN4fnphSd+j26XNmP//srmMyPpA
Zq+DifVNBBOZ7pFpBo8tQlf9ByHxpBF1Ikn4jaxj5mJ5cPyr/9MbzerlLQSckW1s
XETRopBkyd3lfj/pNWH0c8iIhYVzNOKDifdMjjQLMP4Y9dhJ6DFY/TTR9BFkx4ZY
2LIJQn2E5zOYcMuwZmAWA9kGVYvgPXlmKYYTqECtlWaMAyCOxpMLVHsHzUzWHxsZ
s9oWYl2ugKJr7OLTAcwalY6iTpaWcxfjBkKY0j5W20sOqhk//grqt3LWW/fbAk4K
/TRQDtFiydptScupqNBjqahiwM3FRjMjTwTEqtAOPp/pNAdkJ76i5yFpSGdlwDjd
V7GSE5lwaIXrrijQB9PwbEqsmTc2hwqdp1DqW3YIApJAhC/PbkzbzlkaMkb72POe
N9TIN2hKokWAELLKItMvDcWemeLN13/jbHl+QbGZsabcAd8p5DjNnTyfdBRu90CR
VdZpvNqT1UNbfBW9kcswJvOE/EHs6tzQapntv4vmfd8lrs3CJ/HnE2kN0n2XHOQq
ds/4NNS71bD3TupqE7tCiwZcqN36xbxepW2buj1iHWbmYP5KHv0KlbmSidNuJosZ
0rGN5rZSJP4GRAFrTHFZ61lEl3Nfc9xTZ9bcD5ns/F2zq80Do/oSGcVVLUSj3n7g
n67xLWG8uN18HwKc8l9veO1q0nCL2M/a4fsLvZJUGo5XVX1mVb0qmvnJE/A8ruRz
CuJUJUBHfj9d01071Wy+awUivKlTA7Pi0fALaPN+0FNZrgVZpogcDsxRjyCD6Oo+
iVNpUDa8GagaFSbiw70q7L1mqzG92lveCQRgkGi7jjK1nqpMd+CmCAXP/LMvyWEx
JkiXMaWt/zY+0Eb+P5U/zn7qGqIRTNegNF5k7DFz1/XGTPEpU4DDdQJlmvm6NLY2
iWkfAuOUbqwX4YdXOM0iUa2Wv3n0crQ+rFlwToZPMHqj5aGTAgnytyk+ETPOJCHh
te9QOHSGL9AQXj5rI3shHdWfQl6em2KaPpS6+OIguelgA20triQDsEsmQfJO2XSs
dKapGipP51vza4f2QWdhiBi1ncZnRr2uAoWIcC9tZpEbgFAM866gKjaSmUKTurRO
Q6BMOnMrhKNl7U0bTQreKL19i/qUc3WHt/7rETDIRctStN7SNXKwgFySHH2+16l1
Cj5dzl8gyEGLppvO1/yFwKCMYcLubjomj1k+Jw/2U4OypL4hB/cZp+6jyy6DdJmz
ILwNHAUkRkBNOEQAAp85HAYdhM078k0rH002SYymHphu2lbIOHoNNoJoX+x9YRx6
m1UoiW6zSBZRChOGaGLEZl0rZa5tYjTvi5Qmbu0xhBTZukmoDOqwEUQk5KmgbjIc
IQnA1YnoM1/P5OHxZcvrZwJS4xXlVmGJBwvIpUdXY4+nev/v6sARzTNJM1x2V0If
iEdnyOS80+k5zPiwYKADgAhoKHk6nammcwrMeM7qp1M2LSZuLpis/CzRO+4aQiu0
Y9MUXAjgckZevsOKZHwf1rEnywb11agqX6Raf8uWruOofXSFebSWs1HzkcfdM4pY
1R5J+xUgdiT1s/eEcOGXylHUZPOkfQNBYiYcS4xxyR1hQLVFRsjji+nh9KS4U4wk
ZQi7s2N1i7WApWPtuRv4wpuHIFwaVb6SNT5qbmhaVJ7ZPJl9M4zU1V6aMpwtA5H5
VAdJWVki1TDzhXgoPcW2h6wJEIWr0H5zAIDkoNod4D4RhMWDmnVzDyBscopWFGY9
dBq9F9Pe3Gh8zes4eYC7w+J8BXpqknKuAuXhZqgjzLkVz6YicuOBWPJCV3xiVTRy
EsAzmQ5xUFQDE1tQjFhkb+vlMW/jcBz1NPVtynbwbo+nE+E9phcEJH59j2Pm3lCI
oabOPEktVJsV+JOCrB7JSvGxOFq5rIzkinrJjDK8irxekocN+Q8ix5INRm2AERfP
/8/4VhYelIQNxsp/QzmGpf9vkPGzcKGZv0Sltx92fpbM02B0P99ULBUuGyER0OdU
pTOyMRnAl2XC+l5Jj9P0P41oio2Z7tVlCC85OJbmOBiDWfVBNU9TYaMK3fvscply
P8A3OcgeF3t628hfmRa17KBW7lvNwdu8v7nP7U/5Q8scUiwZ7JuE+D45BkJUXjyZ
8RLnedgvB7hdjpuiu0nQmP7ud1wDejHGFMxC5dIarqiRmA4wLlpUOpXue2e2UDMS
uy6wy7bK7twJ3acklg8uV/kruKebom0KmVgsJXtXoAC476OuL6SxrbVUidPB4jYO
2yqNoSZFZkfkrmGMnqFnCuzJq9YO8urAPn9vnx78UmRrvJxHhC44Z0hfqhmMcITO
sVPoVdXKqxFmpzg4d8PfVGhNOGzlfWeAzUxCMsCB03kjom9AEiBNxylHCGhAxjlS
Rsb2W6Wm8zDiaeawdO4lhX9hEEMaZwSMo0LCQ1KDjWlIawWvefopTHg8yTFD0oyK
KmNfjVVPJDG72NCh990FLlwXFxmdb/56KfoJw/UQSzGiU0/YuOM5MSwFEnvcaJ6j
5hOuY78IVN+4bjTxjbe4f2/JV4Khh20n62n8W7nK/7rizq9uZDGY4CaWhno66mlZ
Ou3vSdglDId6S/yxdMhiI4vzpcEMIma0R/A1Rc+VAUQ8jG6N5uysQSh/qIwEwn9F
On5KH+Lg4knWur9t2szVfx3zADW7s5iY9UYicquxe00QY6w+ElXljFu49VfAlILC
g38fiJItxmyHKvekMsbQGFRubd17ZrVx9cfffBey+pTLfmZcx2Aad8Gs0TsjM9lN
Mk05qV7vRhWd+uvDFhC+PbxPhCd3WfFM+dakKguqRxnpW5Y41zjIMAmCZnnxOEue
vzdFFRX9OwVWsVVuVwmBHGKwokcOH7vR79OaeNzs1az4HBGnxvaLvWFq6jPr2vCB
BdKVss624/7bkZ8avPXtgKHV2AyiPFLo7lNHVYjDJ0YftIFNGwEaDcDLH3vG2DUw
/VKxyWeGML87pziC25acVHmsAaPO/MmerNwg2yNWTHMHFmuf4qRp7ZyKWYARFQPY
MyylFy+WEV5uH+vpySxeChgdbJ9B56rpaRZkyJwq6LX3RghFRAp8DSpE5vmXbbI6
Y76wro/55yX74QqwaZTA2V58t3jTrc/3aIDB3eYmoZpH42GU2nF8gss1CnygMW02
ZAzKlUyFHsI9a+RQne71I3dEFsBQrSY00R0xPK8X7OuEqMETeQ3KhepBZnXWYzi7
NOGvSIEulw9p6nrw3LcDrcT5kIfn2OyyrtOR9GbOouQYYPe836ldUVbr2Mm9HAf9
idZGZONpBxWSbnRWOcaUs5Zdmbhg+JGnU2ftN9GFYyTjpd+neVQV8MT27L6VMGN4
C6RIIBIDW5rXNPeKWgeSszq22PCfDWzjO9zmNNGvahsXgIM/YjwZkHzaqqrMf0re
LSUxtnlbowgxoaSrtstkZgZ3dyB76K/A4z5EN5AyiSgMIn9HT6XVsNazwhzq6Fjx
0bmauLaWIHrCYLJjEX7xGjklLgF38O1vQiodaNSaPgStDGjOhYLeOdwsKZ+V9fm7
eRLLeoXfxsLIVOdFjssPj4vQaQ6YtypCqJCvb6lkOHiDAmhYrqTMtdW7mRS96kwK
LmcriOhhJo8ONip7qnRBEsdk1vuIRtc8+Xwp/8xGbiMIxaeD14jcJu0J4hMCstt5
tipF6Sm8p5XEvy8PKYSZufWXY96kvcTt09jQP+24hniI4scgWONktEjEGA9Rk6lv
yINwPWayYSZxBG6iA26fRdZe4ZiG4EEGNssWEQraXw5kyoupjFvppFPUjXKss+Nm
Yfzp/Qoehiufn4nVA8WslVRkZ95G0hOiuYVbwGR45+UwEB/7ij2GvqfOryeZ7Nzm
P7/fX7sgK+p66Iqx6iT0vuKbj0FnxutXkiijy+Y6p0Rj+TEGu/eJos2QLE5ql3/t
Kdv6KWvg0S8bKG8HEjFCXItDcu+Z45JEcRXrhF4hvWVAakFgbvfqEHinoTeESL1d
wZ6guV3/khRGZE6G6W5B8rH5u4m5TaOPi04cc7d2ojFD+D/IAdkvqzom32Kes/lg
3ELhyNBdyqcJnVfOrz7Ko7jDAu8abZGGdLxTH+ioFeJyYDCkkDL/we1oNb5n4ezb
+leJxcWYibckGfRbdDel1ntwOIJDx7OI2BiTJQBlfyboxrz0tBSDj5Nwm8n8EnGa
X5OLBn+9Bi2n25gDR+zmx/fCLSkblUyYT9D6cPGnmzfwehnJbVN2d8HiPcRfTt7N
K2a/UZjsf3qGtUT5Xp4qWTS+xGJcElFNpOQo+8Q7hzh5dpgHZMDj3CNTOS1PZ/Il
bC+3K2XTSPaAWbwoKltTeubsBWmxaR6kKx9HE3YEEZ8TNZhVWuj+64lbw35Rw2Mk
sVXnkAOUxenIQyZD2FE+E+PPhm00QxpnWDRm0ht49EdMbeLu66Pas6t01D6U0xsT
t21TudFYOhDHnhNFlCkXV50UqFjk0I/eBf0yB4bfwGtwS6cWw1xkiD1E0LNnIPSQ
+4OkgXT8NZ8sdjfs/s06hHYFIJNzOG1K1jY22iGLV0J6L3iW+VS3CrVUU05DNvu1
isb6mvkU7O8PIOH23Hx0p7/T292rXiY5kNKGIr4/RbPXC8XagWdfZ9asVon8ar3S
zbyQXuwuMfexJnPmrJPzJeeyY7dDM5y5R8pssWmVZIdf5ejI4QsANpfO66EhAunK
qhyxw+xng1MQ5YkSjwlBNzR6rFAzeKd1kI57B7Phk2ZUzCqKKFs2el4nnEdbq1Mg
OMELGKkXQyCxTvpu5Y1wuB/mf5tQ36PEc9fNaG7M/mqTFHhe+chorYdVrgILMOSW
qKLtr70nud369KY46m72x04sARE9jzAOCGBHG4rm/7tGLPQK4WyWhRyI39V6vDxl
q4+ZrvykoC6CxssWg8gQJgbCXFK9lS86b1ssltKi2sSEhzf8GAs2Xea+/PZgBBOo
Kog3Aon7+j0xZ2zQUyhp8FsZbKNNV0B6k2MLRHzafYQt60h73O4EtkVf7seq7Lua
a+myqpF9fus0r8iK4x60C13bZhYYuJxm5wGHIP1B0vircLZry5sCE2iKFGYQcAic
bjGjUkWylvV7SGGK5VNbT1CeLmy9zT55E9syOHSx3chUVzT7iRYGx2NQ//aiN/YE
MRVDMQTi6RhH39l36L6qPj53HB1LtpkVqJau32XeQU4CUdV6H33J6hs92I2xSxWC
y0xMQTbusXRwhiNE5jJ7gbI/HPunYSSJh9kI+0KZZV6qxrPx7cXEXqOVbBGxU0Qc
Zu8MHCtAG/CsYDj+aIKIYWMU8+cKvseP0eW7gvWNZtwKbL40f1UfKwISQhhuXMS6
4Gz1mpyBnj10k2XaLZmQUFRJhtXLO3+GUG+8ngLVBE4u6s6FS11hUdX1Q6tuTyUG
dN4EyRyRL5i/Ge3YzErQbwPCDMC2tWYWK+30uTS51k6dzaoMxx/Dzlv/Sc5cWbmn
2eh7iaVKjyB7jfUZxqOLEVpwULDko9Emrtjua1wMaIVX8Ob+uBfiSQtTMtKbfw/Y
VPOtZ8Ca4Lh4cGDtKmkr8EnQE/d0ImhdZTjSYIoZKM7Aom8grjIIXI4JcICuIjiY
sEyhqZDLhWJmcLQJJKgEsPIlfa/eblOMweed9hnUIu53mvn5diUKcX9uyUZ6j12M
Ty1pDpNN6qT+HeRBJEwgCATulkzyA76NslYB3+EL5MkuVaTf29WTCUleRnyCDJE9
XPGbOU1M6nHXa5rKqZ2HQ/5E3XngxWhoMENSiLgzn7z7rk7OglWMsN7k9fVBGgMU
A06QzpZnlwLmTSBmVFGhgWrn+CtkqsXhmgugox3er1mxM5Bd0xca2pP8zdiwxAEm
xeojrvSAh2fzcaOp3/kbMekYbHdZWOqQbL3L8SHPcKo9GjX+tR349j0vjtBERiry
jTAbxh8RlVb/x3zgH9GBezd9l9tPCuX1G0vpnrsmez+rzjv5lBX/PUx6MfqVLlIk
+zIFPaA2f0qQIq3RdHvyITcaUfKKasVGkSFrD0rS5zN301CQwmotaXb9k+7XRwIe
mmRbWcbXtmZH6DHTmV+9kPNgtyN9vMq1SA0yUY/JrW+i+sMjLRwr74+8ubO/mYqw
+T7JwzYrW8Ae6gloDyQcm6nnbgM7DUnxZnmUEXCqFYNLUogtR8pk3qiRTMFoa4Q/
L96R/LNOK4CcwxzRUYus4ufa4tt2hwozI9hIQ4/mHtvKY9szqw1FV94XMyC/wh9R
R+z2LQzyUudiuha58+G5qcsMtc5wPgiDXye+kV3bHRxeh6IPv0YawcZKnRsLlfV4
tJK+coHAPKWQ8sTUn7mllZgIz1FHvs2H58wpRWkh/wnoVn6vQ/doO7QI012iKtqe
uxmAcf/vGsBcpVxeKjNu/blI/Errqr+6Ta35dxngSylhs/UDtDZXAuuFxeMx0mlc
jjHLmhdbW2ft2frySVgfdLrO/G9/mv6ujfx/j8c3yRAtAdxUxQxGXbajcqte6FZC
5bJj0w03wmt5RvWZqo6u0x835c794tbw0dXcv1aB3SNUmTEKMW4aESJb7s0FsIH9
tzMtt8HrQ3rPVLE67R4ctcgE+N+JHTVcmzeUfB8rq08=
`pragma protect end_protected
