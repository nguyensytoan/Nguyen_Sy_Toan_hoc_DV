// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:32:00 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mvIyM5tk6+5GHN77UmZ9lsWWwOTvLxtB9HmATEy7rw/RB09kU1wuMSSFvQU7E/KV
cOd2ISiDyRh9CaCTMzDkw8DGdNRX2MC/ZsTm5H0QqWwxpeafQf7LsB6ixgwcrqO4
1h0trWncLfJfOMrTB+zR1Fa/7WMsxUOdiHo90pOuS9w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11696)
SDgvDRS2tzcmE9AL59pTZGFh4jgaM34FFav+PMlB2cTkDS+nnvuG5FX7HOq5wdRm
/xAAM6YV579hFSYjK+8CXOHeBQI7bVnKKu+swBD+Vv62uaN8DnlYOEeVmmm54lVc
sNbO+B6k4XdZKbYcZ3yk1i6VGbMY6PRguAK5AMAmb9/SV0VlwYwd/xIwtrj2oScR
BKfojjhkDBEYDspKt+LyVvPWOIgF0ySjImz/JYLMIA8EQ02MLzs6JzSpMimGxqkP
s9vuh+78na06gW0NHXa7dh5DMbSYTd7fhfsbr4poZNs3OWvMMUlcUUuElh2DrA3F
P2vv1sl4o6l8LWtVvSvEqUTn3arg+zd6zMbERZG6epXsYU9T4H9mxDT9iTy36vIB
7fvF2inAGOyhyJ7WwFHqpgD4D/e3VsoZ+ZDn6A65Z3p70RpNH+wesaz/8fn1N/ZS
zAO56NScyCwxZn0dcbsS6rX0Kj+XZqZNV3rP9Hjqa7SU0VkokaQ0n+QFQt+LckHR
FZeczsVbqHkghG7GGGGRbEr5Ln01nnzH2Q+E6BrSkLidkcL6+Muoyq5osk/iQNSY
52MoI4W3voD8dWOyteI4xRN6nM5mNiV+nfqGH0VCdmy2qnB+fzSsSfZc+JmdDUCz
+6k7Vvytz9VFY9kNT1gpKiINkLDVJd45wnzHUvTSSKDfnf/gqNnyfssPftl/Q1TA
lvlaldh6wPN3+KCwBKFR4cmeJnDUmaidaMarL+SYNGp4cpAqXmSwsB18hBpvkN8H
wwdkbFs/7e8cLMGLfqCKdX2H1dL223FiEf/YHbkrSpy18hL7ZlSsZEGR46s+ATwX
oQVkmz7R3Jgxxd1iJ3+5JMWTKZmDlptw+7PVCEurwdGkaCspWfmw/R8ULa9oNSs+
Tve7W9m4ex9HDEUBBaaQojh9ozdskDxj88LmdesbIVsxzuhDq6X74Tn8wmTjk1CD
W0eOJ3j+2Z5KZNVvRafB0U07nEnKBcMtF//EDKS8bkEtsWwNfJGhRoX/hRvSomEe
AbSXEb7JVDKPEm76Sc5KXMyHw88CSuBgHs+9i90wsvLlGGq1NxKLR2MjUuUx35hm
S6lc1AR9aQ4ZLciKlnWcDYlg4su0qS4akClCz6IQWQplCp1SkFbR+nXC+vBRBm16
r9IGCpAOJ8AsaiVtNnTf4rWu42ddF8cAcM6i5n2iAu2zaZn1Z/s9imHuYSe1OLAg
aek2gDwkE95B2K88v6rv6B+gmFnv5NDI8VJxEmaOxURqtUQEEjFlUR5O/xchBB7P
g4CCHoBKmnnIPtNBjvBlp8AzZroBtciG2I546jmpbDz916rwhsCAXjAxBRpF3FKa
Zkql/VzPeJL1HRgYSkNPTeovofJr4kG5QFJxy72i8LV1OHh3eD6rl0GXk7yGMCD3
W4vjFBU3/GumnJYeD89ZwlUlZMf+AqsfkMQiiM3E2nlAFqWXWSzSWJfxjVHIXB0y
JI03Nu+/Lg3P5juBMZXrbWbPdWIKDws8Eauj+bXbk5Dab2r67J5IOHhC0YtEdsgN
6XCs+5kOE3iQQe5uTUcHfmjCd0U7QrpZhv2UUlSly7UiaJNRYJ5+jagyqCIWsxpC
MzEJ3VDiT9OafVU/YH8nDSWeBwjUSdoKToIEbLkJq62we/QSzPduUxhIl7K55bzh
LKz7sl5zaLvolQnnxFfnXqpkand0VjHprki3q2MzfMTUw0s8SuptHPjFrxtkxZpi
PsW4eoEfsqqTXRqWnJlGvDQATLPr5X1/inN7h3Wu57s9ez4cVKS4zKZvYSx720qt
4/fz7jD0S5sw13VaPzoqB9fK49IeRffH4IxTj8I11cePzJLq2A24YMsvl++uHt7F
L3MzgWk/8nFbPlaPpuVcKKFZOvNrjSSjWgncIP+kB0uq7FBD6RecNpMgmHuGUvQI
WJfB5kcEKOoSJMbPtZ4rSEZV20Gw81qm9jubG26EpmoO5AwaGM7j4dlVP+itTa9F
hXDvNoYBOQShYG0sQ73ZlV4fQ2zUn0A8l9mc/KeRkJZbrxeR8x39lnLPNiEW1aJh
1qByPQnGqoAFowfuxerj8NhOnTyqFAQDo3o38VVfU1THLUcp+oGPTwlOVTF0VOBk
hKMbTCnKRliwcVZS5jHYG+4IJD15At7JZflHwng748M/PcOhRoUe2jfGcU+uzpXa
5RqC8etGgZbJ8RmM2n+f7IX335AWWt+4Jlwa41SwfAoELcf3H0n52gX2neNJIy5R
5RuxYwwtlCPBDlIHZUAf388ittxtfSsq2PWrsKGtET8ExCSxQ4oU5uZMC444heQd
4HRH8P3VTUSADbShajVBo0fH9dgu4Wwy+mAMbqwA6ocWJ+wQ4TbTeIoGezrllrYo
/mgL6RYFEAQpqxuP5/lYLdtojJdEyiLv5z0wuG1jxidNYU/GN5eGr5EhgmMbUDyb
nBgnQENJnbZbh2yo6Id9vhBY72AXx+kiq5RCiF/OcNdxOXWHI4KkGpAmdWOtJb64
VxFaW+JGR/UNNYfIMpZ6WBxQ0jRA2aFdKJcF1CKZuY/FLcqmWE7PU6seB46miQYp
dJaFlvBE9rNMMOrT8Y73KEFBUtMdWDq9lMah32YfQUDKH86uGglrEOy2fVCkXaYQ
FEk68A4SVMlRJmQj3GI+PDrq/FHczVku/VwRvpYvXxVMnUMom5I/j30o8hYSSWly
qwUfVItOq4sUs+OCvWq5vcoL3w0qKg2BvmTJknwfb/dKzpH4CVmoCy4PmEQaIWdl
vqZp5O7xgeA7YYcsVdKpcYiC68OAEt3de4TRoQlM9INfG7OeIQqsaRyVF6KopcWi
L2cOFfrm7R0w1TMpCmljvAjJ1E3pK5unnAFe7nY8ybz5vp7mLaiJyekovjyAv3CU
iskzp7huP/jcMGyxLT9mafKj9kUjPMy/se4Rzvr64gOR71YZ265n48LtsRFYJ88i
FfUi1OoiFRYI+0xnknIfm5C1u3b7Qfq6FS4TKj5gNHqlwq0aE3gbXTIzMwquSd5j
5JMAHedV9Tvm/M65Dpg1RGVtcBLUipKSasfRmEu8J3md+Im0mt83LHJhssDnfN5E
EC0eJDBrfncNzF1E/L7bm6GWptxjZLPaP0TuHKhC9SMxVroauKxVEYJxBrF0EX4a
mUruqGKt5IhJE5tLvx/DcxfP3Q8VrmMIPpCGnSPcK6csjR6r/5LyNoRg+/ZyEpYR
NhWtwwSgDBUg22WMcFu7S7R7b65s2Z6BftSUJZ/FFT+XiGjYZBnUkwjtulT1dFm0
UvFvkpxO7XDLYFgRnRZa5n3xAgLX5exusHqDCWnaXkFWI+iIdFPxGnJCMHE53Q7q
8O57BvbGe9pgylZUfQcHVkqZ24YjCuaR2H0EtfhSt9HCmt8MjwdgkenIHxelhdox
cXjvXVkc34rNA8ZPn5iF2QcbfELZmGlbtfw/5XkdPmzPG0zRkNUwa0+ux/k995pu
3/xHqYTziolhpgjrVl7MoG4ZvdlB3s8785IXG51R7K5ASb7J6VGIDAOTunBs9hMW
LO/sqq1OIHexp+JAmpvoqJ9HaKlkj08JeQrcaqBJv82ryo4/kXCrMP2CoZaDg1S/
NvEqdZm0+tFEpVE4qxbBlYsLxOCxCxKYwsVHwWS+e8GmyImYnixC6oR+YAj801fS
tUVFxLsbwYqa1pzySoGZBth7icbAFa8U/TbRwuNqR8E/QLdlyEezd5dXlhQbBotH
8heBeIU8AjhLKA3fn5aGUO1LWxfPowA5/UHTeGmst8J1ZJbn3ugqBNahD83Y7kkQ
wXEjLfVpWNkZQQnNaFou5NYNkM9BD2Wu2A+aZY5HjNT3eOemwHxwOkNzDlgCbYDB
v0poTFhM6doT60Nx0KzWw+obxE8zLmOeqmnpsdik93HuTjLgZQ1ipp/S6rRmjaZD
b+Qx+C7wfBGoukXniZ9z3s5R6Cs4BsbM0zRrCY0rijCWUXZ+MBpSq3Q79zn1SWKN
4zAmnI43l97GqCH5id2Ju/v7jXiaHVfo+hMLyw4WJMhWOHqZNo1RQ3nTP4FJ8UE7
fOqcUgnuzOFLf05wwWdnnLkk2iiOB3oEyimAshW9rJ02AS3QF7OTi70h3BrJiW0Y
txtv2BDT+hyPr1K/N01zIDBBgln61lb4Xda+RuUkKyT2MzpD8e4A6pyMvrg8274n
rngmYFy9nQ4spsydqNnIP8FVmiX/F6r0X4spWyTvMVkGbldEOvF/H/7Txa9mm7/3
h7hgIs38vs4kap4F8xoEgUPk+2991WVc+rX9VtSanR6fbrvshy3bZINwLWYNBmoa
kMELCb4rByAonuengqN3D6pbCVil4/Idv4e4TLpzEsp9rpPIH9bTq+ls/7z1dvCP
rGfdEX5jsupn3iDKa9FrT/iwwc8reH/EfYigOfVR7egar5mvSnimvdVUhnDb1vLe
MpwN8rj3bSMimegtWzzUIBayjxrnOL2zkheNfjGAQhH2qdd7rr4FnucZDMLF6BhH
I3Z+dgvd9mbJDaCvnqiw7u3FQobsFs2yZ/jDzDZf8d6kuIngCRZfKnWuQsXsBCr/
3lIWzS18YRZGwRN0u1Lu4zr1HxmWwTGTQFAv0U/LjPpPTyeqYVlLElgUiGDSUa+v
K122EA3f0F5X57vxVznyFx28BpM0+a8oi5Ik2k4uiUsNki09ukIssLfxoG9BYSJl
nIOvpPOMgkv7GxqyDfse4Kg86B8Peja+S+8MXRfJyEFBOPYPWXGekHBXkxd+z8Xv
OoR7NPkAm9OYiJfftqk9OJIg3jIY4PYHcMIwrDhgHiWd52a3mRG7HGI3TM7RnHLE
eUH6wmdEJt2KyLKCBhwf3dEm5vJaP1d/2ABBh0aodkZFO+hKoRRlWcgK1nBvsWnE
4zfdhW4U8J4zJA+p0rdtYcmwF3tC+JDWAC/KujdrsEoBvTsRiUumxtYZBXd76Pbc
5B6L5KonoQexI1iornghSlAv2pSfSYGESgtZyaKHkmpuSR4qZq1+PGmvl1RLtO1P
lI3K8Qdve224QRP9GHscIQPUBMYIF849DPwfEW31CF4zwiTDT3XyeIV49sWqlT+4
6wnuy99ME0WkPMrb1PdCpeCMMcHXVCCEcr835iM8Y9/J8Cl545XjgvmCjQchm56H
ClhIiW67+cgHAQ2Kvq6RXwOkSRdgUc0zJjifLflmrQmZqsIOp9adJumH+cDMcG0J
f69FkiFrHPdGiOllwkD5brgiGt3tntyPXQP+wplicoXvVCQ3YWq+O6Py/AiTCN+f
8YqEEamyc6Bh2zKtRaJR0LMz+ID9glQA1qDz8egpOkkkJDzTtpAe4hV1uEni0WSV
uUxxrC1AcWEdwry10nPlJ1/icq+pFzbQrW6b9LUKRFuJWdHNQr/Aiu8SIZq9XzSH
qttZ+ii1MqP4kLOQDbfJEgrxgSY0SjO9jS0mzhtMXWs8Rn7oU35oF+n0k/KhUixN
USanp0CrSfll2pYHblKWQ3roV2yvPVaGrOj4RsvGxiQLUjCH9tcFKpUJhNMbFIrZ
5UgvCt6lXU2KhsF3KgkUM+kWSmTHv8yK1hQ+TjTgEG/2SPx1+SGJcl+oRmQCPWr7
xVYjlj09Ovu8RsaCBIKQqXz/etqGVyu58ROU57dGWBiguu+Lf7ptAG/JifIhVS5X
6BpK75qJtihgFr3kH+Da5+oFUttasXJeeqVji7SxBs8VknuFiY/u9fdoMEluKlgA
QB7Xt1CGSRafHgtKL6Jb3swNnP0IwUromaV0hPIJCdTLtzb4h6g5OhpcLVKy7TkB
+gPu53zUyu8Y7ECc3EWu3LU0uOHmNCQh0v2qudRMoHUwaPPUQksR88sZ8MnWbSJ+
Xcx54KXfKA7fHRn7QsPG6ke0MY47FP+8kbrKXv2tWnOrVycFqsBN7458VE3k/HQd
KfcPmlo4YKLRtSmyz9UpTB7m6ci4GW1yBYOSizJGWyDv1bJ9xGHugbn+WHCemH5f
yu/yUvr2FrVlzEE3AQiA4AYMP9LBwRXH+5sV+DBhYvzyM9FmcUv5Q0O2ZZuDIsiD
yjUTwLaegnyd2xXDmnU83Ra1Cv6uBbxUe4DDFxqt25UnVkidQU1CGOmXkJnjnAxV
ugSvoQeFK6yZaU/+ayIrGuPew4mbNFVMXGOVEcVx98qhcYGC++Um5+Ofjp13KBPb
x3hSNfOB5GSomfs+lTMILpIkslcfxWsy8d2TjmE6MR8Uii3nI3FZJDSRf70LElhb
8LmE+O40Ef9d68SChaO9Tyxo88V3VkMa+7lokNZYQWiZKVsFpNriiF0y8VBvSnLw
Sq2QIRPMhrocbXLwvvhRc0ivp++BS7vLvpJjiBPGXQK2rCL8PsaqYHI631B0w1Xv
+nNLRWi2ixVC8BHqoc40H6Iq4SX89rvGSXIo7YZ0IouxX7TFLOr7ptzg6c5DMMKz
5dKRHuMMyrdpZgtNKieF/7qortJKp576MrQExBf0TjkDIbTWGo5bLQMk5facdxn8
27tlwgldKNssMCkbXPPNKJOHiuPpo0AA0QNJAAS7oesugLw7HNfaTS886P4AHh0V
owDbO3jRiVfNA4fSS/zm4S7VRHCyf//4n1SUSrwryChgI5bLyQXdfxjXjirmKoIm
nHcfTLtCIvHcI71Yr/oy7gdHHHkx0y7VvP37lTy7pL6VGro8ajZR6pPJynrK3AtR
1EzKILz511oLDqyPi9qm8fqLyrBNplr7JHHLzo/lCBNMKSnOTTIE0hL+f4/1tUzs
TaHrtfpkvKHlac3NcImJ4gnWGC1+jcbMRnke3eZJTvo9AWguFMFSHWDeOg0xh91w
+aGTpTODBT/SlK1KPriTXPR1AeBKU3Cdahez8+769wMB14/VYQmCwhNCxDpuFl7T
zCijdeXZRinTekI13r2NMfYUb5YgLv1bFb7zv1OUB2zxpJNPdvuUSaIB0+dvag/q
Ps2zs5pjg0kbUSq6MH8gts2O/o+5bMq325xIBzvv4x7RN96cKj49MEABUsRy7dtx
iknUC2FQWW4eYbbvUIZY+bg3kCUF9P0ZAx3yFJXpfFeyR/lo9nS3cMd5JEpeRSYD
THWDIziI1eN1WoeqA5F44qNqi5JYaGxbPnwWtc5E8d7WCiApa2uUeRahN4g0LmHn
xs96WKH57qGT31W9apj767OVGaic9diPaJNcrJN2UJkQzJ21EfYXbKnwALi73Xke
d5C7VoeeSjb57sEsFwPmUeGlDu/0e+VlvulX93I0YDdhrTBkUEqsQAw/NOu2kZ7D
mBRHrtoKO4PVm9RXNgFFAO+RYoxVxIo4PkVQnCHU0fSSQDOnFZdZImwxleyfnDF6
1c6qiMso+px9F17xpY3ecI66fRmYosLKRSWVH2+3aBN3ww/STyNIjY+Z2bow5fvC
DMa8Q08AeOQkpBSTPvSYINF1sHf/iQCqmRHtbfBoQcv3Me8ZUqD6FoaOnQnCAC/I
g4D4ArahZGKeqaBOf3/jx5zQUu3j4aGkYzgG+sVFBErYbPWZsVlUzEbnbb+K1EK5
9o82W+3llpPxypHjqn705MOglDAa56x061VbkbMmUA3VClkhyCzEPiDKKZ5OoZmW
mXwtvidn0AFkNiH8ghuewH0vGEXO6D+4YeyxWmLuHdw6dgEyzq6HOr1W3/YJGzVK
splMXxdrO02/RFtUgn0jD45nsZdMh8jb0fS5xjgNPq2pGswFfX11gRRiwz+YN89O
s8xF3D5cwUL5ExFwePr7OZJi55bD6PRSPD8DMaS0oDnnQ8mUBJ9jTHLEhAZ0pImx
AbKFTgdRr/aLQuOEG7K79kfeKLDw9dPgzfIYxxWYC8BHPRyx54EKMwv+QekiLN8w
THEtyMk1fQeLBg9TYEy6D4d6pvNH4TGRLOmOsQFyGBDhKaKMZTnZXjd1I7nemq/c
SVLyrEv5tF/cceGtv3e+a6Lz581mEF9itJeM2WXOyuC3PWqCr1EGkSSN8PpOSqjz
LY2jCFF+Z0eW9LIKX6M3i3Rca6IfYFKMXJDmpmsIgEvXoK1nLArDtjMD8o/AZn/S
fq6YeRARp3WaI8GXZym1ot+J8NKSAWB/M+PC6RMlP0mkkmRtnCYGVCN19CODvTeI
gQe9RTSwxagceoqCsED7QyJG4+sKfpc5vzwpCPy94ZL9ZJ/yV7ABr3AC1mNj/uzW
mYsDQoBxupaKJ9MJVf/gvGjDNYcbGcC//Z7n82vqJtLoRarnHcksQBX0fVhlQi7j
ZKBjS9l+AiM+Et++UaW/4O8UqDzJE9I6zd8Qd3ZYlaDADPeWaPvz28vKME1o57iS
rw5L0a1ekRukGY6djBfkrOtyX0zHybKpzXv8tiy1GrX6UnWLyByoOtwk4HpWE1eH
f/uyOrMztN97xVWg8u6uSX6Mb04uWRwJpVrBUf/WFXYa+eO+zsLjzUOV+INuUktb
s9fZMu52oGKjpbDuQC7cwcl5bZbPX/l3J9z8osSh9Mvc/7oN5Tpj8IZ53fqyQXJA
8azm1EoJxs/EExOhQ5tFTM6pOqh/KO6bFE9rIqeVts6JzMwFdhDHRojHAW9Ymv3n
VvewGJfIQ5oEsn2msYhCN8/lBA8LTCEeSIz2BwvCaRQHF/f0VLcKv5v2l6SP6qHS
xKyz66nz8DMBU6J9nVIcAU6GP7O/03dP36i/KhhRvErKnQMLHduhW/EvY5NTVTva
SKwNYYBDoMjAWSmRufGxB/WAgXyfKFVh9Oi6O17UcXLA2ILvysR+rkxf9vnRzcfl
NDFA98DHRU6njoAb2VKsEp8JhFN0JNCTMhtPuC9xO9swQLLBLDRdW5DqNCQGMK6P
HftLNNiXoHroZksuRsmk3ONi77k6VPA2U6sciMKGIWgHl5DCCDtm/UmeSIyXfbGx
cPj9ZRtfSHhNJwfyaw0Xig1ilV4oWIT3x98NMPYbhKse72KXP3ykAnEIZAGqYwTe
tTxpMch0Gn4VwnmhDRXs7Zws/QdGZTACptkzjJVaMKdtGr41DEDoKbIEsAIMZ6Kq
UcIB6LItA3EwrP4+8yAMVsytsUuK1AGnF2JVe/haSBRGX6zRurLRmhC4774vjA4e
9+3X/DfyY9G1VApH9kjqCiHVIOjddIuFxGil8cno+9+XCTw051j4RX26iW51xewh
3RMUI1sDlJF3Mv7docTbSGni4HNhtI/D7+N711rn/1KzhCvRl0B3p38yzriMXvNN
6HBbYC/525MihUYiryWbv4XffAjSTS0HcKSfqzoaIyOD7deCh8iNNKW53g4Cvr4J
IxSqwLbo2WjENSqDx1z87R3giEwvQmcldAyHHt2cYAG8MeL1ofTn0qNxcMqVqz7B
u3+DWjb8jalYgODnF+qarvos24jUZhqiuLrIJESXse0fiykLiw8+ydOxkc7Jb1an
NhwErz3Gi+k12PI/MO1eKIjMtLWEW8EzycGLfJTt0iipUrIlSO0cLVjD5y2JGuBG
iTAyVH3MmOgRq2AutbPjj/elxBQ8TfIaPRvI6Ksy6DKVr4AL/eIEVs+YLgcbGyPe
HqENKKZaO6fKI57OojdIuZCkj3t8hhmKSpMgdy/nHsGR2d6cAbhLaxpoIptl9mCD
dVhFujpUW8Olktp3KHqlGgFR38QnL37+JDxDYALBF9wNowDbmC8+68bvaj9oj2BO
bS1nR0AuyIvpjS1kpMyrOSENzAd8IL5ZqIKfGt001HjDZzi/unwIavDLjdw8pPfq
PkEJYZC2jjwvQ0xSpW0a1wdKigpXqGGvDXflP0nRs0T+6WvNAxFmS8jgGYxESy5I
12Ok0xlPRYtMsPhRW3hNSDj8m+bf3VJnG6rbvW8vVxD8yyKckMQoxudu9dl9BRS/
jrlJWaaW6uz1VhV5JSnVo26+W9rAe1cJ8b/vc0qeSxssiaFuyDuwP0Vs4XYMVgKi
8zyi4XdPANlOTk7qvyaFhsFw7OBKBZKuBMTdGALZSNgT6W2bnhibawjcUinsj4VH
1ddzUaLjQf7/HMlITLYxWlCit099ToYA+r/uvUeY/60qDkCityC8VK6DxFRhr+by
gxFuHxFM2Ib71uYcrNpssH/y9oXy3GjAfGdFMngBDzbv7xvzxGVgyC0ryb52NKN3
P+LXgOfhHFTLFFx8yU3q2Gqk9Q5JV1YRN7Xsesccb6sZu436W1F3wS3/r1WKCkK8
yMUTrIjOOTspEkdrC6iLlgtYH757GmDLhFxCXxmV4EvPZ639zDhaOEfGBDV2X2Gv
jHqx0ncanh0PZ1o39I2YosyzLkcBiZS9wz51wnMvVdC7NHwjD08PX8PTEEQjqiM8
v/s7xfTrtBhEXWLNo/KtOzga1Hl6TaRAcN++FQAHQ+qMT0ZZozr/kdjAwl2FVuaa
gbQlBSmewicmLymUGHefirjio2ZnjCuGCSvYhS9v9h8TOBIw1gKP3DGsk0TPpYhi
+qjSKKLIcrKk1W9WaFpmNHx+NPSu9unbJoR1tO3qt++V3M5dX5Z7qYWYM86/pzJ1
daMiwZCNDoHH7GHsYUL3gaz1Q4nrkxQhMhGJBGCGi6extl+TsJhPqYZgU/sDXW2T
PhutuqsbDXNPWB0NBwUSVO47jz8+f0j4ymNdJQAIV3TTmwtdMsJKsV2sYJnTZZFs
T0VoAwbtYW/EqLYnOfEFVrUu/FbU35b26HYbTP4AKOB3ZJ/ssNCY2RTuqZPeVCiZ
KQ0M+1q9qQM/Qt5hBncZvGtokPbk6JqfIW9EMMS8I7nXoVgTFzfAiVBg+7J+ZCUA
WX/FTSC9r/s4umO/Wg7nrSuPuXsYp6WEf1M//x06pnE2BpW+shQS5aLu/zfXlWuc
4DLRu/35GsicvJuDPjWrvElyfHfjUY/+kpu1o1n3pwL7EzcE7Gm3GBrthFmGfe8R
BvWUcut9p1dXJHsFxq5POGJvB+A3WbqenbeEY4+n8Kq1tNMdsp0mdF72CR00ETle
TGPF5C2YHOGJPH7uS9Fe2gmGnbs+lXILBPBSp2yMeoeEEKV1chLUUHcZlnut7ac1
2dn9dV/rEJz5P09VVtrGo6vr6rP/RSHgem+zhfqBHFRxm8xpfaEDuVKUTai/eI9Q
Kd8/8eMXlS071ItmfUOj0J7ZqswF35DaS0rU59OVjo+xIJ5o3rka4IrWByXKDbBD
QFmVmiouCi1Vx2Ee1MU/74VektKqnITjFHlLTHs7hj6GIy2u2Mt3KFK7lgVgdJV0
FHzdmao6MJ9VPMMAqTk+gNzWnXhbFNrIvHxNQWxHj7rC3SWBUf7fzqlIdyJFwDrh
t/5UAVlG1F9QGxcLV9Py9vinuGp8MXtZTh+NJbl+TMkaTo0Z60LDc+bSVLaWa3Zi
IBDnjf1C7Ti2it4hYoXZxX77CcrFDNlboj+Re/qnRr0JUem+0SIBanV2t+cIx/Rn
RLbvEHjfKz8I2P84uLbVVdqVdhxwOS9zEm4+bqVya3lWRFjXn7/x/YxzBCMpuM3j
yodgVPTXD+3/AT5Yg2ZUxI6f7JhxHdr+cbLpjivI7DidQqKSDH+XmIWpZkmYy7+A
aHav4lKQBBjF8hzaZyEFY3tVcL7i2wRlAUK8ZscZZP7pKCCRKjFMNDTvW1HhEnj0
+MYhPoDik6oU0EB8udWWN2EqWlEm1P9MGcPJWttRcvYbH9LOUl9RjuOHa0tgKApO
vMwDvr6qgRppLJBWCqSAsbbMVtV4zr1L+l+Kasf4vgdZ/MPEUjIeIULnndPV8sgB
cYj5rcTO6WAP7hgc4uZUlB4SZNwgumQIJeb+M8BuU8wVNIkgM8zkUY7kgohCHa7J
CRczIMcXqkr21HyYEvHZb2n0npziT0hqqNGxQAubpVj3zcsovnhLwFAheSKi+WFA
5u9pQwFGEqr+54EtbtKR/PvY7i+jF/c62cmOm+54wIlMcmlPrUuKXyG7/GIEw+ZP
fP6pYXUAlUx2/bvYcYBqYB63OWND+JstFSLvuz72zZaUVaZIGy1ze1myxPXadxCI
pfCdG4FvDZaOROYOxBdNH75bap4/82i0Jf/GwS4pwTaS/dV65M9VEI1qRWt2rSmO
/8DC5xC9fh4bjBTdbfEKnomc6lPvPMk13O21hOURTeBi/ubg3GZulocqnYfwwppK
lJsoEMf6J5AkzFxlmbN0FIlWrvw5ZREhLMVkLr4RRk6Omi6TJRnsmly1QCEYHVyx
/4Ikbc/YSxc5Q0muOxGBugKvl3JdFuX6hGJkyIwFc6gGmgoXeSeJzP/VKiWD+lMB
8UpB9uH6JUadT07l3W2WpOf0xj3vf1VQ90H7vg27H5qdC/mvSnRPiY0oOvmxMcfd
mUY97BJtFVzsDJvK//gUZzTBLqj/1YzmpponGCMMVpvh7NUr/tBZ7U0KR32f2Q13
y9xvXyoQl6t9+AalfDcJBdbtUyBMARpDAxitwN7AN6B0i0+/6dVwtoDuQ4ypGTTk
YNGUUUx3aDaz5TXlc7UJgoFlJgM/z4CUP6TwdmAXoNeiieSEoKeZQanwSb4ACriO
nbJvpnYA9Cmc2ykXW6hDFnJMxm1kwN7V5L34uHqHsi7OsNdFm5mvrJ+znyQAADM6
32S+XGtmkNRPnGba/39j8q1iMW4UgvN9awy40dQHxPvkKQSNt17HgT85KJhi7jux
F0YYaW711f/Tswsd59e0UHSSeXMo3AMiQbHS2irDiEAZiyhL1N+gK/+wsLIGWt86
hgwDUfNm5kzogh2zfXSyqAEbyeTpYw5r27L4qMK2fIOAnNV1Zo6wNVwtD6oPXB6v
jMY6LI0DGhbtueIS//NxguY02Qpp7yoFsJCKC2oCT7pmeS7Eu6paxkCse14hnmlo
2sGhi2n2QEGHQ4GxbrrBfu/ZHAv6VCVa31f35ReJraGXGpC/iMHdENoc4PwbGrrT
sqEsvO3SPIYHylI0I3jrHlo0M32IYpLOZpLeiu91b7xeJtXEFJOadhudGCHtI0Jx
UxoC341r3vnBu2f+2ZCzGEajRfv90vKac+2Ipxn+ONhCOdeEV51Oli8/PkAfSGTg
Gq4RpzgAJFk0WZz7i7ZPe1WH9DLOYMwlmWTXhhryFaWDCABca4mTueJ+GjU7Zhb0
XtZKYTR84CUy3uOZRVWpbD4dGT+UwTUYeRl2ku+XbyBlIDmpyMsCqJP6aMEFHxk4
i4OtOx2qVhPlTO9KVfqa/h5aiOqfK+KavZfY3egxiQdxrOlsr6/q0Z9mB62Wrgqd
XxjEZWJ+fTX0qeQA7pVPNvyFEIYhr/E/Y0L50H6EFMgjhQe5I2DcJmHcdoOzrSj5
PMAd/yo2Q0UHkoWvluoe2FhymNIMI8RXNsaIMyWDixNN28oOf0BKp8t9UlVhr9W3
LyzkU4d5xjcWGuf4QHwJYnusoFLdQu2V/txpFvwRaC/MczIawPZqN70CXLB8XVF9
Tze+iTjcSZ753H7hCY3GaxhIWXTTFWB2VQhA2WPpCynwRcR+/UBDpIuTdSfgtKve
wQ39pzP6y9/HvZkr54evQrjkL0G1So9z46K4INu9jeIU9TklzB2u98ujzzeoiEga
QdX0TAAeFO21vhi3R+FjnXtKICE44DFuTRnKHYCy4OmI4ScFFlYb1aT0zDhcJsRH
AZQZEaenZNeKgBiaKGfTOrCfxLs6ub5DGSYBFzoR2IVr8mz2Un9m+ubqyU6mDKgW
0t+FeOrOGXhzqzZdMeMamfnAxYRytMllniBmqwE9N/iq09NeaSC5hfhR0H4FPAwH
sItCrindvAM5ZWdNB5SfuHa5MH0IGYvPmeyHkOLucCSZaiAr6XiIwEQOFNbjkXO4
61zYj2svmyJEUXDVAV6JhO+EmDPmTnczox+xbWgiS/Bj/XT+ZphAWVrM6r67ysZo
gAQn8sQ3j92nrd6QpTtUbt2lMsAFPmbGEiRszTQS9kcKjvcC1uJvQgkBZB+hEWp9
qT6N4kw6TxSbesmIv3x3A/8+H9xgOeSLAwchuYPGdIPuofBh4DRZPuTECrEy7xTF
3ElIWi9T1adQqcD0yGhnV56bS8K0VrQNtQVKJwqBqK7atQgp0w4g7hujc84tWq81
mOvlD8Z2ugHLlu/zABFi/TAYmXiwvgbNthGauPZIhQ4LsJqT2EF26reYiG5Uv4W2
bAMnfa9SRuyBLY1YCjcHzFFWFinHe5xKwmuXm4aphlc99z1ric94Dg/WZw6Mlgz3
BF+iAmVE4spW5b/XISvPHVEZ3unkCgFh5HBWu+Y/uL3O7xv5j4Rh2uPRpzQzN1WH
X7NoiO7cU878R33atQb3IL3M/eHYj7wNSxLip+8Jln3tUGm5+ncVHr5d8uLvNZW7
F9p6m/Plw+GwuUhuPswia4CsL7Z6ijYuiZzwGKM5nUR8RhozPWhJWB4H5JnmaDZM
Lz4R3xzIOatcwfZQDg3EqaQ368prTx1rTcxpataGQPNZXTuWXKU85J06ciR6DwUh
2I0LkIHvlORqPTpTy2c7iVJJ/DBN/rpnqGH2emdx0SC0vCSAwH0J7+KPUV7DGBWU
UeIRyMUKm+1N4vh1gQjNsES2F1KMIS0LksPb9ELNlSkt/R78J0SUoi83zPA7b8zb
WPLebw2j74rd2HuwSWJ2NTi/64Y2P3NSteA3sRU0xqDwzfuiXZ1fCF9JkNt6OmHU
ZOkJLEYD3OgfEC4Si+H+GJlHpC0J5RaVsakFMUXFF+bTtsE0I/RlMh/TmEW5UTB2
fB73MfDDoYes7kLF5QYDjJ3Qj/oCx+ALIl7bqW1SSQsAZJcaoIc6ue8PxW5o3MoH
Qh74bYcG3478tDdyObfMf48TWCjjEyEaG+s20uYaLrPGcOiMDNe+h2G4OrffGuyr
Dm+aZCYfqt9S7Y6orLauUqO0d195BTHFbNy4fWLtxnaF9Vt34oatRZbhcC6i3M2i
k3V6AdCqdU1CiKJ5+jBsIkIdDIDTqJyBZnjW3DCym7D5v8Wdoc1fW3C8KrKZ4+vn
LwCeOtY9y9nknOHiTrL3RoepALJuI9CTCx06B1bqYS0Bt8T8uGRWfGceMYuSpjOJ
CByvoeSgCeq6ikOygdGZ/YMPG/SxpvKy11rbaHtzVM/aTnyI6H+k5MkKVC9RDHXC
TH6LwZzA5aTN/E6xrDWXFyg7xRhofkF8mxRV3QKMXVcjWGcz4up8vqfkEFrmte02
FwR/4rLQI5gj8wBl2AayOogYBNMY/7lBt2nvD3C1jFI+JQDH5OxIq777DCaQOplB
YNgS4nz3gezz4c6BMbZzFyGEZAEF4nDmM1qwOorIrhO1zvgrniSelSLn/Fyk1pQe
kplfzE03vOUNJtNcDQ4vvmJd2LxkNPDKgESgmFFUBuolWcV8r29GMbc2/wg+kslx
IR7iRW/SWI3IVBBRlU+MD/zwQ0QQADtnnhNmcmEEZ/mZFt5nKQYP2FRK5H0CjmxH
E78ynqie7qZ5vq+mrkdR9ibmZ5HbCEmXhnUZ1yImD9bEMbjgUoV+pQ7+eL8J50Se
+l0E3nEYoK+9cQHgs8PQ+HjGZJM64WIYYBq6fiRQETfjRMYKGBxceUFnGyQc3HN4
/yJwK0HGNfrowZK2AbmpQ82mP6cHZ20RiiZr5nXiO6kvh28Zns855sicGU24QEaj
B1d5hXgqIgSbvjuA3La7+Z7JGdP53ArkQHBxEsTuZGKKwfAz2LtE1t8KeqEdGdZ5
EWK7F+GpheE0LnKGTawxqz67uKY2fCpcIbQB4TTtkWs=
`pragma protect end_protected
