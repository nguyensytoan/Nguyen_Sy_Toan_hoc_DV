// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:32:02 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EJDctAlCODyBBI0MAueqAhKtjk0GOEDl1VsN9HWxNvEJREJfn0ku+ByRKxDcOf0G
WTPtDO6vvysWGN0ik/0pjw2QSghV2l9dA3IEUNai/c1dmimG/w7tJyCzYgvCXQXl
YW5XaQ2ac2n1uC9I0+4kCQym3+K9+MuEQim/8qzeWn8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11472)
nwf/24mPmc5EwJfc4Hpke6kdEY95yQqoni4h5rYnnX5nG4i3pYre1q8yGbq/dR7u
jI6yeubBzHowZZY92ZMJk93Auqrog44ETM3erwvrxMHO8sKxtM69ShDbPvzuMeVi
9/TFD9XHolGn3xpQKSXB2PQPl9wDXgkG8UrkKbC1NY4wSddfhdgwr8/KfVH3ckPG
L3y3TJrKrLF26XgyBLoSyH2EurKWF7amotWuandUZIdRAdcaAP5dKDG/aYTbUEWV
mcFiq0LGlub92ApxqlmxkQYshB3pzKp8am9GrUL85kHjVOk7hivv/YCLxa32RbXT
D9J5bzlLjwbpUYdyP/nubZQsAShtwtAPK1ty19re/5uZ5yTKW2JIZX9eK1e+F77u
xvqrDZwJJ5eUOJ0Yxlh+18J1Qf7X1w5ILZxw00RGusoMjwXXLPvySntUgrYRoC5V
OTeg7ohDvdGxhxPYd5ug1lD4JfspDpZOSVJH2pYZfEAKRv61epXb/Uvg8+MLDTv1
p5Iuq9MwhrBtG28G9s384unCj7l+nT2rU1UuwaBjHdrKzl7w0A53xoQmgumYfb/9
mA+B9/+aZ1IFNNiL8Eoeh7O9V4U7xIG31CBxERH7t7njeHPcoEGytGWj3hX0bWHN
NVMDd/gofCOkxPmKUAFQ7qusUHNzU9SlXy1g6gnxXO7G1ue/MYtu/hQZ1w/ImCtq
Vbt34Oy6Ft7NQnD93EdtnQkDCgA2QTM9essCqAieugSKGLE/UvPO7W4SWAlpicoa
GLOmIQ8v1YCwZA/+xXeR8BUDNzZxzO0Xp0ugNm7mmjgBruEL0x1clbNDHDfYl3z+
C91L+/JZpJ5gDchwSRCAUpUPEmf02ifPKygJtLW61N9cc9tLrOZsA2r4hPvhxKJP
aUjUMF6ETAO6jQ5CIvjOqMIf62MZIvoQZdiSxPsBXFXHf0GoIPuQY1PYhlnL48Ky
UciaKxzwBOirSZ8IqYSgRl6FR4K0wSSrnT4VVL1TBlQsOyJesZQM/e9qpSnk++UZ
fgoTKC5797M/fNOsq9SsREknobaIGW7lbyJOhtrkFeZvcfl0hgw5oG8C+9G+jeth
899v4Z9+zaZHHiL8CzgwX0eg58GADWdJDSdjy5Z1IOPlNJwR7buHKcUAuY2yEOLK
OWfA4hQ5WTUeKirjaPKsorJNOmnQJg9C/EvUEIdkNDWQv9VrnXp2iKwAJ48BK01m
DUKGi2Vt/KZHSRDj5WXG7uMOSebAM2a4kgeQ6mLzbPaiLBJuf2hKUEovIUC8J8PA
9LkBF6ORhATJnPHcCEgA7UwDDzaUDUPPuyRy4fs2eRoBjzZGQFBT4WGbQ82J/fhm
3Wx5Zpptiqat3Ah7b7eO5BjvVrt1r8+RUe594jgc8nzFpd9mKZgvPzIx1/FK4JXL
m9CU5D7hJcMGy+zjsFzK7k45TAg0JYgwQWXjC4/tsw4G6bWuA9HZNrnyo6eQTBQz
nUafBrd4AWaQ9KLDIwSjKOEEyVoPYG7kmTLqCSxjsBACQIbl3i/c63nxhaYp7zpx
VlQt7wEG/JyQk5bz2xMzyUqC274HEZv0Jgn/m1kU1ULTj7tn5BkO3dsuFn28+E8p
eoiX/IqSmHYZoa2/indGPf+TOcU/Nip/hX5wKRm91VPe03EG/TZygNvoPpOq46dJ
svPzkxGlrHpkk57gqSPcQ0+iO1KG/VlKBzxnr+0hNQrlJ50FtJ8AD6n2ffs1ECzF
Ab7S2F2jWhap0Wfl/TaOgkwOnk25q//GMmmdnqfwhxPFZbsSIDwpfmcuA21GcVKi
UWR4WBINidmI5YRL74K9/WAqwd6Dl9sTqMJlz/laJNUBrMHDotgcAtl5U3xqWE5r
p2za2il3cT49kJlPM6nPxIpQKpKM/0/VmX7czL3GcTiN596/FHHaaeASIAx1uKg+
XrUGhaDxDgiVhComDFvtkX80GbfzKkMPi7Zd7MskPAL94MKZsBqgqRafq+kQUxRY
6eeFZAA0JOAxElXWTV/sYDR94phW6QKG5N8LrszmK2bRc6acAs6iihXEMiHnOQA5
fnHeOhCoW6ZWamHvK0fmt4A4NswZNSNELeNJYzySyTjy3bMqRzmPiWw2pNBQwi+N
kZV5PqeAGwUM7buqJl3DES1XfZLmyFDLaeDYCa9D6LG9bBOnTDXtMJdrZJJ1WdiJ
sEyLK7V+SJHmclHsLc8QVZkbdsX6P8tWNiqqsR3AYNalt+y7sweADx8iiP40muCT
NQOe55QFYLGHbkHrPCA8abAZjbp/bT+moAYvUc9hjhx/+OCDfw9EtMA//kmaPvRr
jXihwOJL0OGDiewu3qeWcTbJePJ2FXDFOccLK0m1zW9vBqczHeRvZyEQegfz1p7A
2QbtLlxrjwVjGAyMbULDpaDyYfX3tIl4GBCyLrlUzrPjKeWtcS8EL0QVXmdQqzof
VCBo9miMJ0NJqjyNce+c+Xkb1MrYnzQX/zSs8xIQ0asTMwndqz2QgVkIj+d9ZP/N
2kqc5PK0+rfNBC78bmj/QCmNiX+zwVsDfbh6nSHVtIKpwsgUk5ZUMWgwK+K1G4Sr
pYEr4icOfgzElolnDjrFMAVXdOj0tLkQ9Sy4doE9/ZeTyiZny7m53kZmATAyQAKt
zB1+o9QckwcuxV1DvoxjLU+plHm0St9YlyT34VlRT+2bncdbuqSFQbxEZUk/AMRk
0rhtXTqi9or6wpMCre651U8OBWQuyut3Xm0qMfxB0V3vsSWKXb79V3TYjGDVZ2QM
ph+Zop2NGpbSDbR8mm1EhSDPIlRo8SMjsqt3DOPSTrNMHeG4xnao3AWQZwE8JJUr
4uPyAVUOca/y10m6lZMiBaSY4j6XokqKjfshlZXPXX8IdgXPYzSmfPrEOEXIbgRm
cGZS9vJyxlKYQAgLKGKiUyw/kByOSr7Wh0B/idB/uL6Onjq+SpSHNS/BB/yUp2+/
7N9xy7w+crKocbV32jVN/srQA8g3+3YJS5BxbbCFRQx9skxvDUyPXRTYMuvrR7Ae
ifPXTm6wK3Mjy2oFRTY7K7Dia3jloJw5kk61hDtUyAOsAf4UM1Tzw7cicpMkl2l2
KfWHvhBDFB7GeqIi6x8P9P3/AEhp+PG8zIexBLC4q6LJQWO7uWz/7Fpxe0HPDoFu
4dCUideossDW5BzjXt2liQZPxkNPjc0HAo5MKktAtoS4A8+LnDnLm2N+8TAI/FGt
xfxjlTFAnxrabW8NDtzcT2linm97oltKTmxu13/fBslY6hym5W5dAhyQiOhQcC6V
8LFSZGGTv8G8SzGibaUPrx1gzRcnMXs6iiRwA9yDOhRwC32A83XyxA5/r0pKtoGC
ifNw/aVURyWgmJ61Zm3ADR0PFLXpGASgLLWiNirEQ6NU1NQqIXC9HtNShawJ4hEC
vdNyxQkALNIWdJXhAnyar0gPXkSYPryZQaA6koTljbvaDVI2fgkxK1czqhEIHyOK
G5NpKHpgRGTClF6o5PCc0ziTSTeDeKMGox28GdpMOs57qGBBbJyRLG6Vf7E9BbhY
7u0ExG9egvV5t+QkSVeLZ69P14HcPh0EaXTSUzYeMqcAez6NTDeVuC1G2O1p2+RE
xzwjJo8HUV3p+JEZPIbok7tx87ngqbzDVCW8ILOK1uMqJYUJ7vhG+fBnhn/VGAop
Cwd6V57TBRQJLVlryLvrjOiAL5LQYANPRXsOsLUQ3uZi9ci7TWJnjZHHFeZ4KCKw
bNcU5m0WdaZZBWzwCceNO3C5OJKoVYkMxYuKKywZeOBDHiW/w5xxNV1WVkPPkTps
FPlCClBWt/lb9mCRL2zRqOkbX2N3fTI4PcLb+Fc7pxCyzFZlwQGlvkXujXEwD0rv
iX5UNZ+0dLbNK4BYhpCoGAGrZNkYDIVkg7hxIv3tmLwqqsIo5aWOB5nOJOL4i5UP
0PkLaylwhNUKWqutZhYn9RZKYUm8H9G/TauAQwaWlR7orvlQZ177tliQuhCBGqBi
UWleUvXyeoc+sRpn2/cdQhM8gRfHVVsVut1pnY7Vtyee0FXPLu0GXDVS29fqXeJf
2HOwylcKs7b/6XanCrHT2Q5ElEdeWAyNxEIW4lkitl61yK+cUTYwzTF6EdUvqm5G
xl1hZnue/ySbVuIcyp17Nlc7rAl5ycdkVcU5eOxPWugNKB2z9EB2AZvckQhoJqVd
ci+qan0DNrZkD9LuFDcANEI+p0+fhDolCoiYHsUXF8mtbavk2V68jL4XcRqlMA8O
yoDMLS8ycOzWOyLPn4yNH3L6+HFnOs0rO2vWiFaqDVP6NZwqgFXwzRKDS0Dc/lxW
eHqy3BNdeWcqZ2/MAPLP3JLnyphe3UNwCYYCKgOsohIMZnTdJVG6NkyW5PWF78zP
FDf03pmVkpjQiCDV+ryW3PoUvartoUIgTkln34WbHruaACjbFt8DI6qhcSjqNCet
cUz7DvjoQBXcQzMsEx3qNgIwi/mKIzdsM1t9e6h+b79S8YsKSFhmXwvZvGP7ZTZK
qYXlKWRVKaJI2hl1gu4yU/Ap6WfU+Mel9f0LDH8GJjA471zDDmLt22SMWGa6DFAh
x0trZq1tpp+ilyRC4gRKfuhkW0KGHpPXsDa62aMTZgOizX7AQ5VH1FHgjgC590uD
C5USuhNYNlLnnb5b3jt13H+FZ7v0WweunfUB5ERGMo9H59C4oE2ZN6KTtB+ICZAm
umag3VEz08dSmMFVOd3qSdR716627C9AZRPTgo0/clECuVaDGMsdBSJK7qq8FRLC
tV7IEUzL8if2uh+sqe5EXvBE+EyIPdFjkTMjP+Jb6tx539np/vRuX8GB3TqR9zBN
Wv2to4FyOKq5uRCGH9/IjYUysi+/KLd365YyplUlhIn1CwAd4BRR0OCP0ZSVzErf
+6fky3CFbBi9qECi4T/JmtK6CQrYkb8xRjZw0ckASgXf70nLtPnSsOHz2ihOrLLP
QSd03nyUNHyK7NVACib14MHKa3iPQF/7iYWoOwcaavyIri5Yh8Yg0vnxU28lNiII
xRjcmNHH7JCl+IAKu9Pd9FdpeLj1id9T0n4ghsnh4HABJnz5oU1mLUnaTYaGH2yj
O189em8PZLkPrZ5gUTy+InHdbCkFrHA5TcfP0b42wEjRgiOl0xSgEA8SP1amxpBp
OgqFQptgiZglbyrFfuyEE5e1EKDkRxKlZoGFfXfNycVMY68+nKTqvX3oJtr0Rr3t
Ii5lfNXat89ABvNkWXHB6x6aFNNcM8Io7JNlZF5yhQSSQnPbjwEO3NGEgTyJs4bn
IO4Gt8xPD9eYGqlyXb7QKDohjz7YWZbKTT6ZKBSZ9+3JLd1yaEQKVlsA6OK0DJFf
qi+QW5Orq3IyJEjEr9jZg7GAZ9WNYI6w0AkCOhhSXkg60fkW+7MMllWoip50PAyZ
WkX+Psu2PkdhwoAjOdKcXTd0hdt35gZFF9/w3mBiMBszRLja1Ahbtigsw8hq2dei
PKt1UG0XGm8+GXytGAgOuQBL4TjgbmS48nNd2kf+0Hen7y+UrDXdzrilT/q4JpYA
ClRHf3RZ3K8UHotvxO99H3uajAGwSLY4tnzgsi/WU6ogAjcAHtU703KCI5JjP0Bo
4ycR1OR1ZjMhkQgDNJ3BFiqT16kHwSYf6qVSON/cLFgf5CFMiJYCx3GioNmsi+1G
b2be/rwZlUROKNBa/8zIBrHjh+DxBqU097/QBL5w2J2D6bYMeNWI5J6T4yLY1buf
GUaatNVr2AbyuUZmRWz4W4N36eGmo31YXgCnQXrOxoSEkM52kvYcOVKU6OAnVawq
Z4jtx493K/rmcqTvLZaWN02y54EZjousuxGwn+Knp3O8aXXmL8Mo7DHCdLNcXPaF
bwI6CoOUT7keQ7Z5lE49q9sCIeSVAGSpcn6R6zrSoWPC/LCgohxmB3kTeZW+C+2s
xlWgJPBi/gmNUlr48Eps/ctnOhAsVOnk/3MdqXVT0Ky8tDbhV8UtvFQopknQsFnG
MxAkbWNmyHPuRuhiATw6AFkYMxfLN92hyAq2g7R7S42UHTs0NnpicUkSGpp8sPDx
orOA/8T+7HU+tzj98pgGKQGfFgID8gUqvWIUrZvVT0c+DwhgBPPfwvR+SpWero33
RTPE7YDyHpRUUei+RhzUSy51NEg8n07AxmS4Q2646ER8s6lbP9jHJOpXDeeFgrtV
KcDmoSXzVygYohzRR16pj2xKt5CGHiyZtl+zRYOZ+pRcbaPeYi3yjd6u3S9bGqQj
BPmCJDxKDQNn/3TV1Ct+gqL8KixMthnog8cqKLwC5Ycj4DoIVbwB/zD0C6c4FDMj
07ZXZzaDHVEKqZlRTiBdFuKmm41iEnE3rgLdtvje+VIK0sUDBNfX55erPIds/fvf
jTGm3LvtFIdocqpANRDPmwJWER03o/p8DSq4hMJiwcomuD+wseInZGghbukkJ6jL
4J41JQShrCD0YAyKac5A8ko99MF1+p4g62meoFZ8melwIEYr3auiTC3X8ArWDSkg
rIRVC6kmLH0ieMePUVVzGdEilxAjWrL6EwTSLepojf33ZwhnUZbTMzTdgs59tQ1o
V9nqBFdpTSqj/35nJIp6ys427C4LsgnpAI3zSyrJ9w/vK6ZCDkCZJ+E2kM1hLAmo
IUUc4Nn9DN+8zhm1vd8o+t7YEhfwx111mJH9pyeLtD/is5ldSfo5qGLbU39QZ5tj
J4H5Rfb+R0bWGRevvtUjEM2Zr8+6zu8tLhvnVo2e8AUQrAZxbyGv76LIy5GJgixC
nSoYrUNZ7BHbCbdwpVvY80PCMCiq/3JNJiRgtLmzEGRNNqy+NcDfJ4QJaSGaO8Pl
0MgzmliuGl8T3cQi4242UTBeFQzXUPLHDlQFzEtiFUFZSTKVubIu1frGYZiUbTJV
OhO8TO4WhdnVE9eMY9cZ1eSZIUcSJdurkya7qkiElsDlbVkMqFOhlihzZBo1scl0
AtQ2N39lexWYd+RExsVm240ATb5/NXhU2y2veKUwU+urjagf4iuCU25T/i+Ln/JI
TQdLPoYEdK5R/r9c2P02nbFAV5HpN63OI8P5c3AjSidzaXwJNykbjK/TPqVTZta+
yryHkT8fyHVmG9cnStVDezBUimX3CGkLVqJPVZG2o0+67BW99IDLCq2uxEkDeIIL
OcpyZ6+zJc1LPH8oKp08gBGsGOkm1jJc+5Wpw1uyLtHJrDW22dFwrO/iGlvmUB51
zB0ZQza55qF4Ej1uDaNd2bI2va9O0oRLbu3pMMZZkgbGEzt9D+isULfut6aeCkCC
bLuYpksX6aQRWlhGIYvbeSfYYYPOS9vXyb4/teY30/BfeuVLC2ADoyU0XbFrshca
TqKErexIcFrdqTqab1gOTPr4hszjL51IqS79CFQU1eoG4tTNDcTglF7CsABjQiTE
eyh6Exx/DfwBBwWDHGOwLWkwEtW0sBiiMZ4l1dEQ6zlNg2IbZa56spmFQA9hsOhP
tSfBCnme3CBFrzwT50QHAe0thkkEE0neYmUESvEdy67851mYtFvEMVKiYrmtwuuH
pOi6dosa0BwTWtjmTN0l5YYRUrRi1vOk618GDt+KfL0R5nGyLHEv1DlAlvjChHOZ
/oPijkCqEdJ6HCE/cZDI7JjOcP42zmjoBCt57LLiuWNL1tnWFyLERS8TSc4IaxmR
vR8bnPYEGlyVGWuj2i8L3cG5K5pWmELVBAKBRkpfSg7xzJdvT8Yad8m+/UJHnmDx
nZ9SJRrwU7WZDJoy7a+CqGsrrjW2xKitxBwOI17SUr4OjD6eaWLKeILhstMWup7U
8/04TIJ3Vwdqp3wLHt3yY52OrtxcewlCqM/1Bz7Z2YKIASLee/RAm2gsgrTCnDRx
e1dwkViVPw+C5FjGlXlIX7EGOXmVKNdKYjnDtjrIFEvc66SWimxzZ6KVVFugwqEy
WuyX9AgTpr75c/10lu1ZOk6HBlFWi2dx+mPZ4dhO4P6079kkrv7qpgg9V7D3i03U
si6dbi4zMiApO40EHZIollLZcuRHfrSmdCAsk4nB6ZsD2LJ4mIK/p0tP/dRpPUvL
xx3G5800kkbEKNB+e5t4Hqh/47th5z09sr1CJ6Wzo3xxVSZ1cBLOyqFqBrwDQmAs
sGnfPT2BpqtIdUf020aqbvCcbB7baqojGHkfdzMh/R182XJN/+v4eej+jLgOPDZW
SpBU/Tez/noQ8t/e23bun9U4PvlKrxVXFEExn4H/3aO2yatTB7CKucuv2Qb9r/Wj
euilLA23YYc5ZdjEpLOrttbP6oydks5H3mUBeByABgwQjiiKq9luzpgS2HgItXUS
Cv0mjyLCBc+sIig8wRCqsO0jZdihgYUWZBiFaqFhdO7TWgVEZuQVgiqcKBaFpt1K
E5DeMsGbEHuPKJIzUxnN7GP0RdMLEvvatla1mUlSWbVmkDefVGb1zksin7/v61LE
ZuCzxLs3KyQxezwYRdDGkQJFNA8brt+FZJK0tA68XWowXIQCBalpOyplJe28ykMj
F+9JDmnrCLfhpXuFL/8GgJFHA/rZiHJdxtfjX8XZcb4I3Nwzg3yJnIKw02KbNIpl
quMhssXzfQqa1gKwi/6vArSqkblBvTwoadjuHILPKb6Qvywyitv5Skxp6+cVYlCd
LCM57/YM5SUFByJ1iGjmamOdf5xxwLfZZPsvGtXflf2z/MA9IE8KhsA+AmGFa1PC
evP0wHCliHEej5SKLHEJrIcS032x3lzDLmlutOoLEOMwStAtfQ7R/8swXZudOlgW
7WzBo8nDZAMJAENzkUCK/auehP0uosqR9buJNyJSZgfGOS0rrHqZljozss8hm04N
NdSEK6pzArAmeU8i5IjVy9h9TV57EMymo4j/SAKB/wBaRCPEGolcKeSbMZMe9t52
/TwMExoI1pRDXzovUqqL60w9//NdvxasJzR2sOF236IUOL/1BKIhcbdeQWcyjr+D
rVUg491SamczXNLenyoT+av23TFIPIaA7TBgRAJNyBP7XeuO67hnxQNEO3onvlvt
Q4WReKda706oIsND7tbEBJBhK08g3zyLw0fxfadKMaSIj3zX9SNuyB0JwWxFK+JP
idtA9sT0CkAWTte/XTsY3SG31hQlausySEuayeGE6+AqniYlvXU+LDTO9BVxTVQu
qxFZYG3IlW3GVHQQlwJbWobE9sjUNBI2tR4LSwXb0d6CHvck8UP5ZxTw28ES3+Nj
et3OBd7OvqII5yGZM9ZBX1GUjCsAmsfhboCtmpbV1Y1KRBRB72GZcxBDSpEjujBH
neduC/BHIn0WZrvxtvgmaOWIg+9Gkb2p7lFOU6MlXlSQkkIt4yXTDT6yAXOfox65
ickaUSwOw6v22+CefxM0BmVnktTwotXkv67x7V/A1PRylwFZRogM07Z/rwJWfCww
XB6kADrOH2OAB8dr7lj027zzfecGP3q0Hs+mGU+DLM0Ul+ObjXEe5rCeOC8KRLcF
E+r6D28rmdu0+kzoPTodxHSKnZWL0oltZn3+hNkiDgQXRQtuy386w8Yq/XJ/uFaq
PwXi6kMGSd1tqyx2O5MXb68+ksR3amIixUf/4IxnnYoVq+SlAfJhBJit+mCA9b2e
IB4PzHo1DY7bYnGOs0Qv19UkNg/PX1TR9mHXoNB9yIVDdaNjC9g3qPormt9evkcA
LPCwTm8PjlvTyhJNXXl+rVd4XOLA228G34hRrI+UNm99QigXV8+yZHAaZ+Uibihj
581L1O0KqKFTJGJgu3hKtUI/xugGoJml3Vv34o/oKm9+urWaPu9kOm3VVENnbQ3h
zGZEMl8sOe75PFmjAd8ShHAZlUmAQZUv02hk4EQPb+QUTxaG17Lvssrqsign+Rt5
XgNb+hgHlI7qg2SxDJdfid2XMOhKOd70SzD5G5bife6luOHv9MSdYeS0/dk8MYbX
5n+f7RSwV0pOXUwYcZ3q/pFHreAIyI6Xuv42WfAucGpMRFaUUg5b7KfMaKFl392B
i98htEGJ6GZCnURhnZa2x4pG6FOI9SRD8Lnp4TfpdzjdK95eIjn3kCTM3334ownA
E+un27gg0z6fiicTu/NW5jopQQUPxCVyYM9irld4r0l1YB7YpGSF26D8JV/O5t5E
GSatt9JcG5hTVRABzjWlQM9Vr8SVaRlxNVMgEO9VWsY+LkyR1USNlvJtaOsrpdhv
jhMhO9MS4pIe6h9zn3Oioh/XkJ8qzun0/qks9wazSzvXI70+Wu6+Ooj93hu3ZhAP
6dPF/jyfijWM8T+C0h+Yca45viGEE2uZf4BA6mIXemrlvWMldkgZN58NP6KGOEOL
Ns/p/tpgwTGcRbRcpKbknekCmqmTpFydEMUKICGICHwrBFGYSay/6kZ9rrRhj+32
O6p7HK1nq+445j2WUMkof2tJd4ttWPCkZFo3m7bnkFPCmB8pcJn01FfUrSbWh5/4
Z1MX74F3sMNymc1R8XHNSpvz6cvxfC/G607zmeP9wakFv0plGl2shu0zbxhMm9gk
lwoo3jnwNJdpXA/EAjVtx6viiPI9ObVr0B+XWCw+OlGr4PZcmu3Lt6yKx3ySxfbI
aCQLd07askiyhSr8ikGUGrpTHeszs4XRrXfLnRW9GtJuVXvGmDh/sKvaM/4cU1+b
Op6BVDLaHgsI240PuXg8Hs4o/ImCvKN7AovD3pLEGBqv03uZYG0PkcOZm0OeoXbH
Be+VGhNHdzWbTNYUUuOH48LsOOY1ThqKnUVgcsxzatdTsHzFVutIVUyo0GgKo5sU
bfGNM64v/NzB9M94FhDAtvAEvcr7r9X3h3bvP7idEw4iso6hLQcmg9TnxielxG1o
WQeMbpgTTvUj6Inhq6N2q9uMExiHTEcsuemzjnmiwKssW6UeKLrWlQVDQkAhAJub
7pNZ8wifJXtwx7aeI6rd+gSFC8mBlnLNCOsCBuGVEJN3mEmQBJHt+O/jFW4KhUZu
DZy6TStXt+ratjiVVlhi4LufSWZn2c6YmdDcRhBQaqRo04NIn9suIRG40nbsAM7J
t4jqkkPG+YwHyUIK5FNNMP9ydd+rYotntxsHpmWZndxC2tMbD/0DB4LYgjyyQokU
HwWe7SBdLOkDPZXlWmYz9GiaiZDpH8ZGZQmCX3rPHgNKeErg0r/mzE26qmhV8Av4
K5m8U6ZR+3zYTc4Bzxz0RB13uH/vq2D3s4scDm4aIQLtbapQ0xzZQ8ixWgMmjU1X
iTxe54798sMXMDDvGuta6uL8LtQyQObfFEADatFjCxK45t/0F3/5AxZ9U14PJA6B
NzkYQS5s7CHe9k3VKYnrgKUhHUjOSvnaDlqhFvPBmgfGt+VjaFT9dLwTEW/tusQA
u6JEHv7xruFSf5w+KJ6gu1OxaOvRFzQC6xBA1bDSxUIHTPq5VlTNMija5CBGPVvx
a58eoov8qO9XYLRCzIin7sCwE9cG9P2QcbPlDGZDrGWH3CJOBwZc95/RdlrbCgM9
G0ZKMT0KBGBUl8lmdUGYIZrn0jucBcc4kkDsLOUgp86hMC3J61a8DSmnpCZHXJs5
E0Qs8NdG0WvHTvorRvQNOkmG3RcwHXAX9v6jlKlwKJhF7llOkJzzJXYX4KIicD60
DXhdfpZparbRwhpyuDlBnWkZeL5KE++2+KQuAeuqCUtNS/rBzEQfdCfCtL4v5xnb
f1zX08IUhQwriBVgH8dN0Hju+RuJAlvOzWsPN+zRFtBGXCo4CLptLsXqXUYC/Qvy
VzfiXN2bD7hLRGUzakjeV2mluY9Ns3vf+Ex3qxSTsPEQhHOo12fVuFKXIjfP9V8T
64LCk3nrKTIE+A+cISnB3tg6p/7P8nx9eJQmq/5MBODfGRB8RfnMh7cTvQcuK/0+
xWoG2PIo17+XmGl6nOUCqVkincUpbQsrJWz3kuLzTS/yKqlZgi60tcsGm7n5gheK
eMybi7BxIxxPAWquPBBVgVDaZu7Wd1W2vcwYCfGkVKmh4XKzT7K11FaIJnIHc0td
EhqBHXBnE3pLwX5PDygGxNLH6qtX7y1LA7kUx2KduklgyFXJ+5y9X7mnEH8bk75q
lTH+JME55V2clPubC1Gs3pgoecrq6X040smvkkH/PErhQmG4LZVdQNMhZ65T286P
kWy3dq0E4/DohCAX8NNnp3yavLm9SgqDv/2B5dyp5eKd5FVaj/U8xFIaJEHnf/pb
H/mAk7JWLqAZEuvAxKliKMLLg3q0cQle0VD3E01Ws2mIL2OaERr/vL4eeYf/SJpj
XQAM/LnW1ZtY8iEiMBtnPByjvRcbb/kxnSArwuWkpAjrqQEH/J3I3SdJjGyivWiG
pE7sShM1ikYV98wL5RG1cPowJ29GSOarTHNzrJ5CB5GdP+W1XfW6EYWjvsChumaR
bT3Io0lthL1mnymODyRDlnJxf1WdKjzzC8wi4kMU8JFzvmAESEiHRskhF0lBBk8g
LJX7cPLX4bk4YdSOh4sovBX+KoczjQ+JLbeFipVnljcqf6x0nqE+soVNXvMF/1/i
XLtlxM0u1zMUUziWtzyOgBDYaylosgwLPfE4NSHgJ6RZtTTma1oo5843FhJ+nnLC
t0dU9G/jwXO4ASn9lc/TnAvRvoLn8VhxriE20ILsoY44Opbub56kKuJhvEsE1Gvr
8gjltHunTKUx3asD3LwzMEBpXitjv0pHalJdKgivx7efUd8DAYoN02B4F5mwgB62
D7gf3gs6Y7xqpoa6vOCIo1ze9nwKQ90yXtFbN/L2+uvyBvR694/ZwaqfzQ+VacoU
Ed7KkI6VsChFFLTCAn1BSvSJZfIGDQQAj0jfflFTiUu3d5ZXMthHPB3QcPgPQtSf
s4BAbPE786vgdn5Ij6Dt+WyYadagatZ9gLqfayUORt7NS3dBAxWmAYk6i9kjDhlK
K+nNo++jC8WREDviwHrBFrugzLlIacxrf05hAPk8D+AfZWQgo1IGVgy3mz6MadOT
tgXkBdgj8LxsIPxqYFBz12KtFPp0lWMMaie8Ng9ceFVFJtLb+I67d3QugYO76jYF
UHwUbiWewH6doVOgugXFR6UztRNj7sZLGPntmPrKSvja/1RarKgFbO4LPfei4W3E
691BgMzKx5S60be0gNKufZceozRwq4oZoXed9FOzHWCfeK5MdqVJh2e5g+khaHuF
O4wPCmY54EyfOmUTCTW+Zbvw8qlvH7Rrk2IL6nJNkN4PT2xiWz2ke1BMixtjLnJU
J9nabXssdErLXz+UxOWRw4nFTM2zMZrnQW1MGOoVSdRGAN4TBtqVUCPEHy7S7ff5
n30L3WKlcXT3St/5nf9i91sIdiy1kiYDFl18rzwVZhS/LeyjaUhpBeCbXnE6EaRQ
IYMz7k/FDa5atD4XUuM//o9/SK0HOttK83Y7fqAkHhOVj+HY4KeWIWB0Vu6ny4QX
OtOUHbCQO0oDbnIEVAkAATMB56VwlaqoUylCLNU0tzhJACC+OGuaAwiYQytIErsE
ylUVVHjUJUufmJngvwc5jmPGwFDWOCimzCMSge4xv7eI0p3AeqbT4/gvaP1CFNa8
NWinW/FMwYamek+dpeDP+5cZVTQNZjWzBotUHVIRUVweWl4ZuNX1gQQaLV0j6r9/
fQ0jjIO4Hz4vUhL8RIBOCLEQoVWU4qIr7O9dUSh60pvDZ3879lv0ojYEJT4LI4Vj
LlXa4y1Vf5STx/kbj6QlUjyOiEzLRJm1/2sXYxq189pDQEctzoTpDMFSR7pF6Tot
62qJoBpPUsotnJ8Luvf/46QE4zaOx7Jd7mzZA/qHvSf1oEnOTl6UG4SR9eZRo9zg
7C4gwhpNjNPdS1BTOdDP843e/Kj/sInRZU5idg4wUgmvzhqXVTZ3Hho+F/ZZAw6N
hsxhCSJ92EU/VzRAKeXh73JOS8KYeYsbtKtQ+fHV9kS+hwNwKRX3b2iKwxw+c2gm
Mwe91sDBY8WLapHmdMbIqgvtbW3dkYdryw7JYWYbZ1mnvLbex7n0cjFtk1jTBmGa
x/u6FU50NAnToMw7vImFTRw4Lm4TyfSWUTlQHy1gactBJaxe58OiDceGs/HNohLl
vty3gEi72THKaZqBmluYtGLM7tNuVDk5jq0zfQQQcoqtN5BiqAD9MQWt3yqUHVW8
2YKxwA67c9igaJyWW7katbDBw43/Z+odrJ8fKKegbxRCl4mHfCF4MFjVES1Pf7of
t9YC8CkGdMfML56ftBrg5thEZSq+AiRhGqpBfl7+KDB5AZ4C3CiGgp8LqyQR4tuX
BeLJNB4rkUVK7eC/mqkZLZ0xaXO1lJTgB6SJw/k+LENiUJqfMbJbseycshjfd3cK
kDLZ1XX9WxsiMFxMmnEHOLrBMGV8fcLfQYCbNhiMvkxpCDdnIdGLN+YHCMP60mkL
2QvfHNoN3L8xaNP6Z+Eh+DlkFkZyVXQulFUr1vcqWlKxKYCGJ4BjuI611nVbWW+/
s6mZI1MYTHdRyiSRzD3BlYUecNSb17Sjz/NIjajfvOXFeaSpZQCX3gUggPaeCUZR
GI6F0Wjlbo4k8Gkv/HdK4ObAOhWeYcIsGb4RpdWQweCs5W7VnpheVib6aNwKyveL
zGKWfng5bK66PnO9XmorRptzHOw/PvQIDMULEnbCjLlCTaFRjwbmlfRtcwDInt0+
zmyb0oq6c9x85LcMT9lYuR/ZrZVUn4wBIlnvz/kQTJEuKzkv22GyGfdA9cU/1M5v
MWDWsLUNihSO+Z5caooPhPnJdeR6E1WcmA+UFeMf2gMves+O1/P5LNLVgGJvKW/C
tKDqj31FWZ7oiq8Lv26rUxDSzFGdWjdr3UiPiqkmPoxjt8GgLdXHLLBtW9qsiRWH
tyMdeKMlEQfivweqBeJlSLWLP1a1WC01AqAGJAdxXZdrWs9kjG859jmopLASXxNR
pIMu50LWABLXJzwTf82eFJDpqnGrTY4OkON0YNp8E7iQoLZjDQt2reiKLXwu+uHK
XfovduDjDDyVevuH6MuMBVZqRvuQtBEn0k2IoHG1ATBPyCsWF02MBVp5VlxFfE7y
ooP0ASG/NiwfhPR1CDKfHaEx8OTNsnSTa4BuGZP+KMeDxC6/0X+XL2pnThRouPmR
XMZH4qa3CVw/AFL4Ho/zUvy1UZWJVlbshf46iajAf0BFaxPZmR2w06H3PX7tdCO+
zBdkgRwD4k6LUM+MFt1CckitoIJHteqWLrk6h0bMq2wtq9Vo+7d0nxRDKd8TMh1N
1GvJnvNRtyn2tw8xmhpqVeAJ5sPSoNgC2/Qi2BK9JzAonsU1fvUaj5oQ8kteaMUS
2393N8W4JExxrFY91nxeuB65f9Xi3DVYxVzXuy+pmKmG4O5OrP2jL0T+TxxbuBMu
WB6wYO8FUq5iRkUiLxGZJbFQilRJo7YGRM1JJNAGWmfEwd/TIBWgkLE5E2Fv51iw
`pragma protect end_protected
