// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
YMxzBbvAu8AuxC4IiweZv14euzswyEmtg8CRSZo8IIT5mXt5ZpP9DPL695g80Krj80RSVw50EWFM
NwrGGURl135rSVaJz//fCHN3RxfvUROJgKAz9clMez6piHAVrCc22gwld6vTU5Ty2hBH6rgMQlGB
qiEzuCd0agnf6OE/wSx6AuxrkqotJp/HXIwzWhGAsM7Bjsbdwq/Q+R9d9AnTT8THvGo9uJJlXD93
6iLjpOj6k68X2fACrgD7pidX3vUTS6lASNjAW2QIns5+eA9eJoXfx4927f92WBFNNkJMcUP1xqwS
W2o+VkN8XpZKPPps2DR312WDXICg1njy0+VEpw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11392)
iEO7ANb13SfWzBZC2A6fg9J8NzALcoalt8L1LK5Z6XxGhxOUz6pdjoJLX3c2NKpNQZm0z+K2/IE2
GKlLUhshS0UtmRNp4NtJQ3bdwNqfkHF4GHKqhCnb3EvAKlXA6QSkMdFs8/+Wx983VMV9CYyu3L6l
a5qptlncZtNNbrObST+60WrJytxJ3RSgG7j4axRhFI57tkSW5DLuNhrXdM1cx1i8JXzauCjfpdK+
slIcGEwlYJGTwQ3+V19ZzhqyoUDtlhExuZo8fhKaqdku5DMyQ1ogQwLlsl/BWImfsJUUvqxJazjw
BY7zqb/q23c9jKMTEDblov2brnaziEHnIpuyqqPDRuBce5xdE03onym2uLEAJgUJiU6l+r2zTe+z
mT1C5I9oOxKB7MF5JWDvoPLFP/MCc10cBWZWgNsSDaEjhtVGROv0cbuZvnZt2v3rcy5rw4ovBiNC
w9zXFfCnxJhRew7luTaoX4QcP0OZwL2fT+sUgn5lyndMsJ3b1jmRB81sJsvPc0fouskEz8aq+TJy
JacoiogasLT9rjd+6dBvwz9oK3ekj3CPkn7+JRdtY6q6ohGFDkV27aMrjRiO1tqWjU9zcV/Zd6Hf
0zfdM3IqHVUA0w5hDeGI7SrXT8kXa8WcBtvp0Tf+h6vqDKpBNsVDZmLfVx7xKuIkFVq2/fI1b2IM
ZhyOyTmu6OTLTtbRBuAxI4GF/bp5QEotgKHm1zec7HvYa01Yk8gMgmvEao7Lj7/gyuTS0YepZK2F
OFPkr8r5e9sP902fOy4BHcBR0ohX5ks8rbiz29l1GHIjyGEsEzBgoq6sjyk4wZRtT0AP+uXbIlDS
bnDgnxEZlWW1F9WjO4UsUaAi5M+zlG5x9mDngLxl5faCtWosjlQRQvJ4Sm2LnUEMHQ13R8AyQKWu
4ITexN/t2iRNCExviUj2a+HfE+Azb3sqNhXeM5pCi3r/2C9wIrCBLPqn89M0AvqRRUy/Khl1nB5i
3C7p37el4b0IWW9Yw8hUnimCm8kKiMBk8SSbz52c0bukMgSGsOHd2a9fRjiLpWyPuxhOCNexXuMN
OUCbryFE0SJVpPqKN+VMd3/8ijzKu+XRCaVKNerTjmCvvffRsl10Id6ks57LjlZV3fXG2pL/6hcK
terJ/vc42gD43/ELFW7aLnuOX6TXYor9GesnE+8jpk0RqLZFI1t3zD6J2g8UqH/bCc/iU+GdegGU
k8McpeFp1lLSsYQ+rZNbX/OgdJE5TRgdN1BTkNEVRsHPyB1d4SvvNzn+9RohmpN14RKKuvvV7Zzd
eqtHACXbaF8VNrP/yp3/m25IEylcCB/8Q9j8q5KaUT7PdkqfWW4bOIAA2xFkwnB+Lq7RmCFkuZ1x
lH8cBUB5B0NpM2FgBYQqba9pzg9UqjgKQAavt9cvIz6i6DCuYxTqQ24fc862gjA0fr20E/nnYHDO
ZkMZB9lQLeV9BNC5QkDWtuBMry3rpYyzM1IhDhP5sQNihDpSqpCjc15HcL5Yyc6wlYYjlT3EY+Qf
vZxqEPPuzuZU8bCScKBZcMMC1nyfKSEhWvqRxQ1zC4IUuNyasAAeAJrExJG8LP4+FLoBIjLNFD+R
e+RH/W8mO9o8a/Mvezkzm42lDEKyWXdT/kRzo93q1vPYy5icTEx718UhJwOX3gUyIZVXPI0VmqMi
ut+TePkNuWXTdndT9oyTJomL1X7xdH4uXZS7HSEtF00K3GR1z8MpqkzJdV5sYtMfxzoFWmku3Bvf
v2h2ZBYECvbHmNHtsmvcJjlUHzAEWPn9Nplcb8N3izyBjl1UTykqBYw1GgisU99Si2DSF3uCJQjC
WyuxVTSQRhO48WC4kSoZ19N8agEWJ7DueSNe3BhS6vlP4DbW6am36Yval5qTg8gbC2klwTgQwt6S
tJfxwRJUsD2AZBX2mvKizQRA15EgBaIefyZCHA7CoMGsrH1Yg2+8QrK/lgEYWTOeIWoDybehpC5g
TCG9rW+LkldDgr7SmlB4iP/QkKyUzTTC3Q0eOV4lq0TgteBg7CSAR4jvY0uTt/I+SZkYUtk/IHv3
EDaq2GbdcGheDvnEBv1kKbTzaBsaQ+uLxfr2ksE5krDtA745CoXdY+eH3H/ClYZQ9rQzyA2R5rYz
g9UVs3ZGLCCulc/F3pqAw0ravded3bUpJLN6RF6OdjU+X1DxuE+ZikcmtM2QOmCSvZ2ECEBNMvOI
UMy4hjDakFHHcUqbJ2gaHeMsS1aYucq8E4uB4Zg4Hh9yw6Aao9RX5iahUM9OdF8MPahNmmKYVgqJ
+k6n71l9x2zN+uvyZnGEUGbWfKsfXWv+97EwtAiEnCk6TZ/PYdFyiiH71xGgER8LQ+s01/7OPtvc
dfqAu08pepAbr+Yht15VoccVz8ZATMxAJExmjKbojjY+adTLkBV9L34WUjGQXyxqehDjf2GcQPZT
uLPKvlED3sc0T24HL6tTDV5HnNu8zUf2oXE8O87VkYsEAHOZDLWkrlwo5x6ppqTSeIBz3iLtYKKP
uIoPL0+le0YnxaeU16Dbyp8dPsHlcWjpVrlTNkw5Se2Hi+RF2KT/CVBXyVyr5UZcJx222iGuQDfF
LCuYHEGd/NAZLaK6qFENSjhYHK1qRGatGdQgWAmGnPAQRkhiNecjz+K3pEWLuAeyXP6bxWKud072
iPtyAO9l7tlD2ObGH3Kv/ZVlWCNrG1pK3+INQKumdthNvssJKSJD0nyKqHVUdBhPEmtv7+QCS/F6
h4+Y4+83x08BzovbkvM1S0mjXbrUSNnevuk6kXP5u4M4uxJd2JgUYUhGNp7OgF9eA3M/Cu6VsqiW
WD4uj3xEDngxsMnui8WmRF3xBM02YCmV+8TJW4gO5Bms25XmztOW/EXuEKgjTDT+sROY6Yeog71o
LKBn5l8BaigGwfq+jKEE3LvLHmeYBChJbctxxPtd3reUQ9NBvOhefL/vX8MWTusEbW4DIF1f1hKY
fTpn6972vRADp4DHBK1EabbV7OFxqqpefIzgATFgll9TmBMDPqV8hzPRvzjv+Yy5yVtcKCJ1baDO
a3vnvEV2HhXO94LVjonYMNS8kKe99/3uOeLAhf2pXDj2aNgQUGI62VtTv+qUdA0XPJNElNLN/wkW
FlMCGpHRJV1/tXSqYbYp5jkrXzRDKZMjcQBvNqrnZRuwsc/BXqGMfv+RZ9toXgXvxbXS8By6//pW
4aQMmjPrv/m2uN3QtXgOaTRszsnEmVOrfP83p0v3A19Mk2/gQju9t1ron96kHJkbP76WCIQUalf5
L3y+H11mkE91LB73B2NcBxdy3VZ3BKRTrPAjUOhlyyxvh+T27Nn5FrTGdSDIUCE+jR0VSOIDooxI
cmq9c3YG4QGLM2HCV1rPmXHSBezGaKUmzDDp4AVeEJS8GaWfPFxpiEJD+xSWVoyMeprCeCh1qXkg
WIPD8t69Rq7ZZnLfEJqj52y++xSpuVbk3pcmLwpWNZD+gkstkO9BEADNM4UKRT/1a8ex9hLWhU5+
RyqDwZ0ZsgX+as+cTLhHBft+e7HUNRCYvnWqPnQyB0C4A0YH/JhsNQBpLjXW9yvPS8LBrElmz+Uk
chHquFqxVbpB29u8Vg7BmGNhftOZgSsSkUG//6ZC97wFr6ghDr3wLUD1GFVmYMaZyMFgIfV6XMYs
WdFd2/YtqycColZIvumqpGYpTtS7t9JnkuW65YU+/yTHrrCyD6hP3eQNsJ01XXJvUfpTIPyTVbOh
h/mx7Hw1mQ4ZbTsu1U7+/2GJ2ZcaOrzp1KT+QWqLbo4htDR9ciKJz6e5JAKwaniilRXMHauK+Tan
ydyzqqfQ6Ux7B2FweQEvOjD+zDNXo3aRd0gfwevA1S1NJNiUz+79IUGutdvYOcG3kc0jXFAd+oxX
ULS4A232NK7g3PvgF3bUnmUYUpaLrFMvVSpPkoLEQPDjTXj7ru/fQdmVcvCX7spOabP12T2IhkPT
ddbgBkiqkr8j3zg+Yyv2fo66bDZ7Gu9qH1Aa2sNcUp1sjvI1rNLHRnO3e5uZB1suYK/TJSeXXlxP
xSs93yTddJqY4Ken2u7QiiQNN2H//yEGkDn691teW8DlnaQMPoE9nejyx2TjbKdEOytKQBzF+fbi
i4rD3ltxdGVTgNNZRWCen1ZgFsh5RO8RMtgPg9wyPCEpZpfMnt8bGPl+W3TmWYPVIq0y2CuP3sBo
yqgYRx2OKpZUJCI3gOFfXQuxdG721aDszl44CbBhnKODcLsTw0xf3jEcmI2B0fuKmpDz0MAnMpJY
LZutil58mpGXnLP0RxrzWeq4lmUXniXrggKBWKUepfQGg2UDPT3EIj4bqynbDhU9eMiO/Zdt4dLh
+Qon050b/IGs9Y83HyPBJeQvepqcqproTNuXxrg1Lv2NcI7IfejPtg9maLWcy0IGjF/2OyixRF+f
hX7RTzCwg5tzkJ8CNFwZLUh0FzVgmEEExW0fv80NivJqQN4EzNn50OvWDpCCRaf9KSOt7W9b2dxS
mVVTPB8aPojqDcJ1+kgJ7xxo3qj0GczNi/S/jhxTFsDVfQ1zhCEiwVPjXnMeWuGPr/4rKRFwq/6F
8gDdEWaJpKabM1UPeM19Hl250bmauFT4bW2vhCdUj7MMt1kKH4CU2uNv7cEWDduvmWMCpOoaHvw3
hVwev8+BHVEb007MCr0aOM0rxRISLEJEBaSEQRoXLZDH0ac8Ye4vQek4gOTLoK/Q760T3GUOxQEg
qUI5uEcCf3CFQIGKaTSeaKBz9+Uhwj2Rz1Kqn0KgfvYFJqPURd8b+a/qIviwkHvYGVyKWECd+1eJ
Le8wbm/4t48bbT1ncED7VHDIJQX4c5DgnC/fFZ6BfyCN2PgC44mf4+ak0Rdqn1n3AY9ujwX7zNtF
m4gQNIjgGgRxhaY759tVInPFZ94vvXdUC2ksyr0/7/NKAT3iknUaWcaDYyK16drqJzjTOwnVGF7w
EyvULQ3FSNieRBoq55kqml4vSdGsEScZvlFp1JdRmdsR1c3csSuryMXYqOXRh2j90Ox3n5IYj6Bg
4CHXuIvydSHSz/G8citTDAi/Kz2G3xrT1WreuYxDMk65sCEOPH5cYtlIEW1C77bh5ILoiV6Hrbdj
z5LJyKZ7mM5gIAvIBNxz/WenjVt4dZILiwSkIbwMJhRzesHk+Jx6z4019C5lNlron3aEQxGd34wO
h1YpEz/L76x9Ll/e7uOJFV+WBvDkePxYfFRAczsTg7610lEd91J6Q5hnodWLCdAafR0myRrNwWz+
3q8CkvNviYlsgpURjuPaeVo3FDjZfPjMPHW6liCkS+g4+aGLq0lfjRy/WgTFG4PeWTNVXcw7qHKO
z3mlYDyRdwFVRwf6jyrc52kCLWke4tGafCGDSpC2R9TqlmAOEQhdlpZ4xaEw8bgLCmyoUdWGWzOU
RnwH7nf0SSUc2gwl6bXOH4ggHg1eTLy7p4b4Iy/cePIhKuT7mo9he5OhnBbRU8RQcznoiPG2grjE
6Z1Hkb119KqTPJVXOBGkDpNehG6KfsCf7xrWFt+ziZ/eG8ExlCX7QR22K3kOpN4I7vW634vdGnji
xjWpgWbK2h5WMVcfxOhHHjAt/4bdaH9rUMXscjouSyjPE0XKsxSbCPB0LT4fEUlSBwFgAOSMwpib
NsctERSfq9jB7IAbzzy0okS7ycjhvbbKH7MFUym7yqX3lbJeSZAFcpb3PQdFCO6lhnzQJJLDOFlQ
u481L2/FtyPscDIV1nhOVFzPdh1eGHm2CVGmm/gITgob6MVSCIVqJO+yOL/NHbAHhCNVlKDlGC/W
MgRNdh5/OYNOhMjDLFdNDcowfcJFdwNpJ6foUBFRXhn/wzWCgJqkysbEZLRtjsg5fuyTVd2Jf2ky
i3zqq/Kf/8H9kbbkkHSrV3FqXnVXsrnST8OE5gLFst6UtZtLs5c/jBpujPd1jLPKWG8iqytlwfBH
VCuvOqTKzsqK+e1Oue3NoMDN6hO5KEbOkjvkFX347U2GgL2axCYjHNCLNfBZ1n1tN2iNiqsI3Wuw
tZwumeKcPvkWv92+7MhBUBGjYwSXVcDjXO8PqYvcKsnAj7ONKhxRq8bv0Aa31xbK6fIloboTi1O9
YQaSc+dw5RvGhoN1zEJwJvAcgjUXVrEu85YWlbHzLOPfKMKKhBMozfoC9xzyHUNUZGpLCcgVjCAl
oeFlR0dx79iePM0tJZQ+FIR+MuRmIEeYSQJsUwxusH7s4Su0rDvXRHoUwmZ3Lm3+zCRKGLF0cQ9T
nx5NorI2h8lyfPAbPBGLtG9jXR8SojW/SnvcwsX27BuOHUH5o1cLLatSiFDOVx4kl9PLUcHVlh63
TAVF274D2X7xJZ5I4di+BVsdj55zDawf1jJuVy2s+sHEa7BY9mFFtaplMx64BUeI+HOKbQRo4/9x
vhsqt0OyLxHYevBYroRvHywyAEkyP++9Fj+hgrakiqnx9ka+yc+INs1A0S2teQQqb8csGT8HRtR2
bo1f18nMD7JPSC2LxIEq3L0w+1Iu8Ky58ucRHKywvavQ0WtC+10hLuTEl0PZf2Ev3kFrUuppO0+E
6V+Bqd8fJcQNTOaOM1idi7l2KeTVb2sK5sqgkGmXc+tCS2QCSezHh7CfV3nfPrYiR8sntkv99K39
wrQBwBc9axqLqAWFfj0L7pPsOprHG97mdnoGRGzzqTzMe46poa+KIl/I7r+73Vfbka6Z8vPAET5Q
+PuddLr5bsdfhWiJca8ZX/PC09tpxsq8nKgEOMs5E6Vx0YcK6/OSNLKTRJjkNAx9OVdV1ZhfW7JO
cJVkzVBTaTV0m/8+m8GaEBWGAStG8IcNA4ktEnPs3AKFOaG8cQmJv78A/9Y/e+hbPtUKP/TfNUMp
+yKmEuo7SOpQYsoK+wviYxTjDt28ROydsSXVrP17LhsAZs5drdjgtJg8fGvFZVK53kGPrVe1dNUK
jiyE9ML3CCVoGBU+CRl9UITfDMPIuVQiP+VPcVIP8Trz9hz4tA8Hun5sghtxVDbRN1q9Zw59X0NY
6B7N1Wsk1DpnLXhA7Hv6sbiY/Q1DbUn/9LR+7MjQvw2TjpHZQZstTN5nq1cxjj90xW0tn0wlnXIL
0vI6O9g0swVcN+1SQkmvQOfT0EDdaDFSQohjCpIBpUORYlXHMfuGHXpmlxhKdDYXs91B9Z/F0sJv
Jw9LEgsEtBY9Qwq3ecpYM3gr06dllIha2Sj/4lF6bNbKx+U6SWty7xKdQ7sJqGoAHscAzZLuNv0Z
oGmd6Shy1qJfUg7hNnuYtX+KKAJgYtoflHzj+X1OlZuk4it3jrFk+Ys9lZignCnI3PwgC6lXvpKU
QdRiasK4gVtbgvcjuFoJLnkgserEwpg4SgKvvkkhPxIIRraCD6zDNbEU8+dn/Sv/cYldR53GWNeE
cxwjyRaTNCITvy7Tgnw7/q6Xf9WSXBjxzDwodYyqLNX+oCoYDdMmU584n3v2RYgY2TyPIGX/VUOi
cw4sfjxKKsHHKyqnxLndM243qsIFBPfJG8Ltpond+wFAb3mK8Q3UXXWBt+ZWq1zTXxWTXJVkcS4/
/yDxwQMVJKYqY88Wh0yjQA/aPjHJpZhSqKNTwVTTLVEeBQbjTc9U2orwlLeH28Nh28nFi8z2rIlE
O1LoqLn3F3dqKc3/FXPlIE1sgjXcl7N7GG674zVtQnQLYhd4qhXemzkt/ZObn3S2Rq+FJyXo98Tj
4x8SUdHa/htZPtrRGGU22EHHiu8bSRj8bl8NwHPk5Outaml7jYt5Xa1gBt+pLPzT0Frfql1TJlWq
6XPflrnQ1bo1y4+e3Klo4Q69dyv6MgdGdfomocVS/qxnqFWOy/6HwO2WmsntIxRZh7vj8JLcpbPc
JTu8UOO6imOZIl09zoP/aLhUponkp1Hzz0zjwuMESmxIBccG4QGEtV6vuRgmuBIoxPWJpAXmMb1h
m5HQdJe/UzVWNeLbJggAEvPpcbdp5G6o5Cl68yE7KK9tD8b0wldYshcSmyBtKVPL9VzdzCG70ezu
XxTJhv0dgPY2m/ufsKxsOMSBpxlGQSvFhrEOIuFJteyuUZ/4EWVWqsFDaPRQB1FVjZji02sV5fsE
aYGxZs7fwo/q+l9laWtOb77XoUi29+AEEncyw7G3N3rF7HT0oMtGkYw1qOnbJ60S4/E/RPDfIKyp
NDGwvM0996R7uFJ799PrQL7Nrb4jlrZd9uYSFEtE+kUd3eZXvBG/IiqH5P5ejcyI6WORhrnwCIEg
FXnVuLcB0JE7l3/N+6LNH0g/Jqt0mi1TASjlNJFbVo5BffX+8+gIdOaiSftbRx2u8ApyS6t6Q8iJ
wU5P6HIrEHX+V3BVsZBqfYFeBX2A3rjVeC9efval/jB4vNALxAipp21C13u449iWoc2oGUeYdjiD
H59SReIL0FOoVoLz9ph/sJ9BZLplza7yx+d7F9HzQEnm0ct/lG6ZI4UdgVqrtGvxESIFblkg2aCm
u1KvRRLI68QKZOGg5+Ta4PsJL3bYydFRNaw2THXJJsdte4/g9vZaBsHQqFrUC94s+c5TKi5WEXc7
uVusOqRiNUwVoWT0/OcIoBzpt23ikWO0IX5DsgdODAw2/WkR62M/NrRBfqqRs4hIy4u3gShqYcxo
FpwQQc8i1d+sbxB4+yzO4cS6r/8eX9E9XwWWL/mWT7fOQLz+IuOY/MjjwgJgAxME4KqHGCF074bT
gpAQSTxx3iHEo8VdYzlgGQz2wT962A9ZhNTYm6s/QnD7Ugln3J0zbkIIxATn9KRhnBSkqdD6Lkqj
jxSZXbavbof7NVQFYFL6cBpQ7j9qY8m2i4JK5c2IfWDKzkFKboJqRdv0WOw0oewTn9rVuzvAlrmz
65yoCF3b4XAMZodqz9s8kd9yG77lajgvrJdB5w0GMIFCAvBK1SuxPFdmSnRw00jhC/81hVP1XkzM
ZsP0zflmDFR3Ecba5inLvfILLDZNT8mzYhE7PQs1J81ru26np9bDv0Jayqrk+NjJXyzsYbQLu9MJ
altThAHQmcmevK1nH1ch7e0rJnUFDrLSEdkLGPSiwSQUl81upmGF1dImKA8mU7a2xcmxo3EyQfAM
g8c3aUytBknL9oAKNgQ9K1DooOrTaqItZP42QOAhBGcZ/lP792cY0LDK+yTVJzMnN8fCarqXGy0W
0uL6zxqI1AwfsAv3aaPc/uUrFzt03V15Mr3nCbtMu6PsfZknz6xvpQzRGinZdggEuF7F0LfDnLV+
qffDzgXzqr2vwqd1+oyiCdoIneOMCIYkfc1FsufWqJJd1OhsagkGKE4cUN0uZojjEHkuI0GkbBUb
c7WLeOAAhEQnfWZiiPnwRtyAGS2QSwysSBrvyJXw+/wSKFMqFVg2yx8z6ZhJElpxbL3R765X4tKH
4G/PpmBdqD0X4qsAiQsFS8w9Hm406XiYK/EkSbjBt57fu/ICctSdcdXV/c6ucMtnZb4FWi+kBIT9
rRjrrFwDQuDoBYf7xZRuoXtTLPX/ro6fOPixuE6Ro6PEKkiLBGS8ArwJ5Hf242yzdjHi9/gkhIlh
qC9BaWRvY9rIVOhLpxgfVWBrKeA9yas/jPSy4uDv4hG4s/fJANp31qlU6gZEUHM3K4v4H6Jz9WML
7gArpZUyJ1XQju8/f9er14aVRZClfgeOUGBCG5fekyae7dzaC/Q+jCA+Ffrs2DvnfktfzxOIHr55
u1fREhzWv24q/VZTlO2KhM35JV4HN+Qr1th0AGENS4z9QNZOjDZmSfkyRkx+3JZXIqojOe2sPbKF
WSn88Sk5biQiMKUKXhxXtlZ5ny2rbwk2SPwrnAqNIx5hjBqRSoRxeohfa0atkTvvnI4e5y/pOSLe
RfbEyAqPnzv/aUjhxL5A8tmm9Hx6tLJn7UVcW5P8bkVL2E7wORJ/RRmuRF5oEiYrn4U3mE+tjwzQ
SVLpjv1VxLRmQznWGiabXlX9hhpoGl/y6GCZ0GjI8BFxmTkotCVhPN2QW6SuerAPkK+nCMwzEOeN
1bPyiyq1hnVGOsIz7vSPWH5rfCPB1WLG7eA2hdw4m/qA4KYsIuuot2L5ek+NBGhkQ22GNkJlfWOu
02ZKtCI6SpSQA0ub6b+Zv0DOj2pE4uiJynAYVPGmAZc/yocud+xa1YK+hBsqqJO4K+MZv66glh7D
a27Jmukus/JNvF3wSzVOC4N+8b/Sw9S9rof3pAI2I9pBfbtOy9MzS4c2L2flhhmA0I875+tgJsss
XL2A4noymLEI6zHzfezrhcXAMMvuBL6Fdgw+ZyzfgNAgxKwQnermF1sIS65q4gc6H/855pebPQLs
0wyAfSPoKOwrvyWiJn9wTWNEfwZFAbBGEeqVLfN0F9hjhexf3TDrx/cU8Xgvy2jma4HT0l/7Cl9N
et23Ve9C6wgeUE1QnK5/Ww8s9I5lDl7sx+hKTMz4VO3KSvpNhlR6EdE0hSnd7aXqnlVJfd/4k5Z/
8zMBNqjLiC+WUt5FP3vAApqGiyq19MdRsNYxEAmN3iEOV9lIUFdjFklMveYyG2eu/VAJA/Rydh87
7z54EICDIcARgIhbishBJzd4HqtwziI/tl8gDR8XV5H0XsXJfHjhMAf0eCnrx/M3NIm5AtEU2mSa
+hcZEd3RYK/9neBxP0mKtgy5vFy/GOTgSytUN1qqu49c9ZtknaiDhNbRGEmF1pY0GBe/dO4UO1/v
5VEB96MBBJN3IqWmvkNTadRRWILutOceu/95U5xgPTXOOfFYt5VHhGEJ1uMYQHZmtj3ZQXEQ8TgY
SyzW5QSBKCM54cawBDh0VrKJPzPaFJDfh3c2wQq1bT8jmqPBW4+oMNurtK1dncOFy9s/lVLTcPCw
O9tFsU7o2LI0XHZznGa5yFqZjjW201KnaOhyO3iT5QUwkJYB1q9httPkKABAPiQeX5+8rtg9OG1J
ifRHNcA/M6KEvzR39FqY7x/zBv8Nvuez8p8vyiDdLN65lR203eSYankdMu+73emv98Rsqut963Tk
fBL369BcDy4bwJKFZcBE4LlL0MlySxVtXETgz4gca/55O8a5sxXGq/VZEnHK7FyznXcMvun8Edg+
eKgcxYF2QdxWcpj5ohegJD5OTBtWd0Pma7KJriOXgkB2b92jRlHAntkw3K+sjKZaouZrWIICbhvt
o5sFUyhgV2uMRu0DP+c8BUC3HuELw52ZqLxBzBim1n5v0zvTvhobaxRLfkDm/lvkrNJt7hAhSnJv
5Oj6cCqM8r20RcqXMJTz10bswlIko8B2JizdXEZ9okMKqmF/fqKSmK9D1nCkdtfmSZ+8k65lP0W6
b9y5TvOoFKsVeFmWNp0LfwR2t+Y/JtMrLRzcloyJI4xi6kBJoJ6h6b0h5GkiMBjLoJdYVGJcjsgq
cc2nH+W5Sx/04yrMo2bQ6qhccEuYCv4k6crX26u1Ca0fcCNwHj8S0H7Uk/T/UsQZ7pQx9yEm3p9y
hExI4zaZtUTHQSyUMAZ78+AdL6X2O3Ooj2T/MvFoY0kyD4IY4UxXcBwRCEYruUwvEzwPYMwlgCpz
6t/aB1JWm6bhPTQt4E+IMsAWp6xepGARUTntpVLxygDboOwdi7gSRId5WNUNyyAfayD6yM9k5q1q
p+4Iz9Fu8EpqlqVUALGBEZU/2enaqWEsBFcy6U0QN+NBLOUIDIGMTQ6COB0MIc4GtTvyG2iSREVs
suclMjcC1qKKwFjBp/5I0GmMDccmBukU+i0V6TblqneXWz2kHhCWbUSx5Rluam8vj+27mtSzEoFF
vQMoRUEf5AsKd3xAu/d/18RovhzvqnfCzP2uEPUzad87ohqBZCjqqbcFf4MlbMA8Ho6ZCbtoVqFb
tVdp0lKc5udeejvx0TtwSksQSQN3E8vYgB9cZz12OJdfnJSx+n2IFYC2xHkg17tPxEatuPwOK2oa
I9BUPOBpQFck2MqpkyQI+51od9f2qpVx3lkEdZbJEWFFKP/aRyCQgZru6NR366pH1T7XRDCguhwD
8YdYGSc2wgvajiUuLekASVuf+E2/XKVRCWUWiq0GHt/d29RvcTAMbb3B9R4hevhtv5BLnM9MTMAM
vEJdZZFuC2Jhk12A/x5UzMg0Fp8f632YxD61LGbxeBLMm//a0il2kiYvu2KYMomfNsG/pjIA//th
B2ugpOjM1xcWQ/J9j4ZQskAmSd4rCUFmzpTe7dB8iwBsXtsXcz6CgvqwpYjM93A4B9BVjV2qVyCo
34421lhdkh/GiIfiTepN9t1eXrxqIxXL63/gBUF1+iotx45d51XXQ6LtV+OujvakM0PSZN1NJTbs
Xa8VMRMITP528373Uf9KU8ZB3vfbHhMN9SsnG2Eva6zWu7ZK1hnuXHnlXWGlJbpXUk7SFmQYjHWZ
toBKvinSsyo2aw7O4Xu1Pad+qmlDO025IERqdD+2eGl+1uhadjoSCxaF5zW5KQRlsMuuQrA9SeEu
gOXBlbfgIY82YSQvqGtTPuJ9uOhUMv/q3sa2ih07+mmcB6NtTeEt9Y85YxXghwGCiPYwD12CzIGi
qqUIPLNXf7lvDfVxCRCA0PO/How/tzhNu49CXS+VhUmGLZkvk+seoa3q4M5t8fuMf+YF0+m6z+G1
fdyO+dCxKyo0vhtHBclCeX36gmXEdfcvg3YMZBuyRVBiqA6JBt7MbmybDfq2A8LkyzsCfCjrpo2t
VDyrF7P2D0mn+z9l5UrSCHBMW/I/fKAhH7x/ZfvkSe9RkVqnBkksN+pHCEIu3iA4L+wkcpEuhDNv
iYXFJhuAINF/kcwT+GWhmdOLpok/TxIsO1BSWEogPSLB6PYVip4FuWAn5aoy8DkEVgnvPt9UauqW
PpzvqepN6ZidXpnBO6DiIBVuzAUAuzrVXDJ0f1Hi8F+8boyZBiBPOIoVORky7HyGTQeoYgl7NnkH
bNUSxlw/eKBkJ/27yg/PUANjAI8qhirEUqfko/dUTl/FdFG9+EHxjts9n70RoPmbeLZrzk2sU1Jj
CtzsPZWnD/SFLihoGSUvC6ta29i4YgaNy8iF8IK0A77Q0NWzCGSi4X1QHRl+F+ENwpMws3xiflfu
W6mYbvUR1QLrFHjOEsYwvwzJ8CQyR73gefRx7NQOv1JLF7vuT1PS5iDGld6+x17jkFlQkFS/wKnr
KBx75hOBJDST2OAni8b04d5CRGVJdQNULGJheLKDoUWmOXRKLkF69RtgYoJV4UPcSauSiBPK1+yP
PkTIHrOVO7HDTzulAWX8sT4D6FjYjK1DCkwuCpGDKzUJhwM1ovlFsvQD0GZhlaThy/7QyGtL237Y
eEMAbGeZmXYcUDN1SKfW+2AB+ebAr5YU1OuHSiJdCd6Icf6iTk0GJ0VHkgqRZ2ddRvDD96Nmrxnh
4ZkEm2rOslXewtFOkA7J8ssbb8kNy37j8kYMsJ5ZjimHhQV79XV3/T1FvYl2EPKSnKdTqhrkNDCT
BkQQ9WjdIOWcbPzycviulLfWCGB1bQfz+My11c2VXINPe6j/10Z2Fh6D5z9kPgcoDB5DEtqh9Pof
P0nGVoQIxNFvyHHqcWOfzcU1HMzYM9nXr0b1sQH6K/1YtfaSzecEgh1Axaw2JVwmF99wsHjXteyC
+jWuCPe2zysnBRQnq5m1TClKHKQv+ti+WK0euXUpTfjR7JR7PitLxVRqJt9LGmfEFSkkN+vcEtYK
+zqaV+j9blKPd0K6uy1TN4LAj3p3fvps7gx8EoSXgGhXlFN14F8cUTd9AhvPlEmxzlA/EBM2IWbt
akRU8xxiCeIc5XxI9V8uQXR0TK1Wv87S7/oaVlhwMSqGVYQD5aKbM8aU7a306ou9uye0/FSMzzld
eFMWbRib0jEPWCaRoC/AzY7yKJEfn0idNTPCpSy9x17qo42oasPZQhumOsCyOCBIJHgcpVi3AY49
aWuSS9lfEPHGEmMMALdfy6+3eqE9lvsFfpYywT3my8nzd2LR1nRna3OGmWjK4X715G7HdNp8ZvRN
RwK5VvNZ3/1QXBaLSBYYdFQqk+zdciqE0joxhATgqNtQFLJTV/amqQCHa6cguS9Oc2ZILpfKMMXn
nvrsQLIpZuJxviRhfHDBjaF1YV+Ld9rZwCLd9TsVnBhl9AnB0oZLyvlekAlsGcIzurnut9RaWEGq
jvprDC/pcA9fZWLY0Ts4+8Wxrf3kHlWVhnxV1D6Qs13x47xynUOv/cg+4v8UGWYNuTJX8J7UbPuJ
uxLzUhuvTs2APx3Fip/aPDVSi4wwB9DlJBKWKcBF09RLwpHqGU2JyZyxRjcslcgjbT1KbiosqRb9
QNe+36sZOwZD6n3hhVNSYjf/5DYqIz3aIMSwIpz8811C0vJjikB0lXapTxWEqS6vctXPTCrkOwzM
dHo+znAacOxzFvu4zpTDSIskjJpPoznIeJB/PDXwmMrfm+1ly2Lr6S50HBMY+os9HgdV5OSqQJTG
btjmVzKfuTFZqc1dm67cgZWqJ6uga+WJluJAC6VTzcq6JMGKZpHukyJK3t0r0S91neWIQB7ctGDr
11iJmLjZ2aFXxmCuahIbrb6pte6MC+tbooSRLILVcgD55vnkaqu8JoEhmoEo0OkobIjBDRa8yPsK
JulQ12Ca80TRrqyaiH1OkEZO7ucOwHRtMTb0ZxhdtMy94rDYDGxxnmTaNz/wmHjJTVPHRnkC/dGG
o2of0Z4cj3ZA38PNN4q0Byzwe7PelhtzJvISXkz9RUgvvRNzz9gwwBtmwOaZC8lmOt4vOEGq6pHQ
jQwE0iHuVqLFjhIRTRLi28tdFF2w/bVxev544+YIGTjvL1ZelQ42kt2KT6u0Wp/1ZmROzjcNjjdJ
M2B+S5kewu2ThQTDveam95tECHDn5abXvBZgmBYrotMZ14gqnUxXtcwZ0qlwCzPlaWw+lf2YN9+G
jjvr8wnviBwFMorKrvGeVT8/Sb+LwDv8IFR+culhxkM86qysTShMhkJTQDcNxS6EoLypLCJJn4P2
HArRTxniSu2z+rf9dfehbWPYHUme0ZfrGGScQDub6nq1rBJTkwDX/MUeOZkKRh5Yjs0FdUCQ13K5
H4yIHKX5YApoMvnw5iiAiYxSypclgtwGr532DDRSHCNyL1gAf+9/x4XMB7pcK/N0XB6qrDwWZz+4
/Bf60Sppq+52sDkFiEyhAGZzWfr7qySZF0c9WZ2FngXLP4KhHS91pMfsHEhifTZv6H75GhiHkhQa
EkTMPFThwUneiioIMUc2ZdoGGwNi1GA5exRrILRSAdzrvk0Z2h2Dl1C4CVJ8+5bF9Q==
`pragma protect end_protected
