// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
X5mpyvyiep6ON4ABU/m3xWLhqk5/FJVsuG7FblQwCHNVxiH+GQmpPSFWlSkBckHQVBjFXy9jP1wy
QJ17jK2pCM5/lcEElp97bE8QWi0i0lXIH0aG1DXzWjS5s/qtKKUWpsNtkj5fH95Sx8zLaz/HEKj0
O2FguSty/3O0xNAYU5l9WNSilGOrGIy1L0wXD1ZE9xfeM50AOuvzv7Fl8ndkWxX88uCkW1DJI1LQ
SJEkg94K4bdg7LSZ7lvbItAdlHNGBVZFdze8t3zD36rpS3PovJZ1G4aKEXduJTtrdU8E27CxgKzy
RsNzpWRpX8y4uugzAXMGok4T+mUylv/IM0ZCxw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 17360)
diS4R5ZGNG9qD7uPYj/4w+JgmkBNKVVssK49L1lVbVK5lropQVqb6jaqYsbmVQPCJQpSQRd8J20k
2rcA8l/V1i2ZDZJiKYa6O2L/XVgVgOeoIpw42ckDi1k73YQODtrMPaVrsX8zJWrzMnmGeaXVkAJc
fUtDoZiLnwu3iXitNWb3AH7H5wrgKBzqs4lAmqtNbSSkO8SsFCDSnR4ZzQKrzqMtNJX/CUaRO++i
bE+Ic/neenv3TVbtYrNxQUL6B/LR3mzsL0K8rWQZROHRQx73nknvex86QyFRRvhz3vu6xYF5Twch
uvVVqdOb59K6ADWPbtugztddlb3qKr0V3dVDlChVuGSAV+oXwl/KD+sLK/Ck5LuUUm4FXChMY2ib
FWtqRdgHGj4BqmQWBH+/koetkTetjBcKCTtqLOA6ylDVCzjJJu3GKS8lvHqOn5SK7bG0SOQnz5wN
2Uw26ueiJ7rokPcjv6yVNmMN/uVGWx5JrK6bTMcEAo7/zYXA0yaKfFQYjQDcDAl34h6RSpimjAwQ
6WZtBbWVLZIYaTXNlsM9PEgmil+eX/Y0z6RJciYlMVm1wqOIMlQnw6r2C22IelVnQavt81lhroql
RVpbFigbJmhcTZUOgb4M6oCB+iK2novBEfkxdrff+OgXEQiKZ+/vLk6mVvjkwYD1PAKF9KAbWTh8
5sPURU9MOfJ0howrIrzrGtS1PWCGdTnb49SEjZzPBl16221Sa4hsB/kYmvLbPJYwHZoSDjWp5nes
79hHl5kSydKy6AplARwyW54axiO6rXqAs8f16+o2MTwyjlaUaBxFWvHfamKt0penCm/vOmQG2YM1
B24JPUuFP7vO6JXmCjNdsDvNzOnTbb+crU3JuOBMw3Cak3rqNgZHg+XiN112hyu8hg5Qu4eCh9Db
x2iehGXWYBvBPETNrjvR1vndPQ9UcUekmayjCYpnaib70TFYay6uIXZbGGe4P3qPu6rFZRuzUERr
T/yCVFMEApsw1hPlOZjKlvHAae1dgrCgWj7IBqMpnryGXCXyMQkVCt9n0uIv5bD2vBItyxw6Gcit
hNUSTd9F3a25hi79EpqGvNKERdHNcrGFqouQw4c1/PRQ9teiDTO+bVAX74edKH2NTPjCKWp7Tddu
3JKaPjIun3YSj+CjTnKimd7SNkoyi+tqFj2JYiF3OHWkcbgfD0vkvY63XuWKBosiG5oJqJWlVTW0
Gu9nJiOpDYVT2W8RZzk5qW+7UJ0BBulNzjPbJLiBOjSYGrqWjzjDWvcDhX5c+mO6RU4DSppj7l5R
KVaOhLHqu3TI388Yl4cNPvpp0698DyjCHFqZ5JWY34K+sZeJJsX4Mdpare3I4xLtAxzj+0f58sCN
P+Bxl1nje1aUMy3wmg4KvJeAoViROYa+LuUHkgLBWZ7rp0DYXUhLEYz6Zn96pq3XpeAtYSNSOXRM
au6EUMwHHfzaW3ylkr9C89v5lSlZagmGWKBU4dNnxshpT3ebs0BjIN3P2sLg1oMvxzha043vQz9Q
MxRqL1XLDcPeRizDyZdn5RTJnkT+uRNeEYADVPAqAmgml5Z+FOeFFnxPmzEM6j2pmCanxL1DNv6P
IRazmJVw8KJSvg3KS1DtwCks53gEAchybyvY9wAp3xcdpZE/CHcw9To06G6y8GHRwhrT4SMW0zh5
3F2XcPXNhcF60J8vSDCkzXnrrwog4Ggswy64cuYm6CAe+Wk3igxVMOvlX0Bn0igB9iP6Uz40ttw7
MX++4ogYaPQYQjKuR0ZZ4mTX99NbOvQCWPrUT/E0rLqsBhntpMkuhKagA4JrS3nkJx/3OH11vVIK
5iw8wRd0nKEX38p07nF3GDOVvSfTomCgi+FjbyhlxANh3UQOe1Q67F28ficX9JNElVmPczI9Ezhg
wwj4Db9Vb4cucSHsTgjwXzJI532lDERhAHK982aZTsZQ26el9jnqH3t2KjDLWAkIZ4Pe4mTnKOO5
jewcOU6z6JI1NM2qD+P7TxJ1C6L2Vv5lFpgf+FaX1VQ3cQHQVpqLg8pOlKcJ6BfmMbPHuMK1+Ahj
MnFViRy3EZonAxdlLKiBWVn/y8MouLtW5CkYhcGvkpqdSQKqeUVf3GGGfTmKiuXY1NiVxW/e0sjF
LMhBhezcAydmGuXoAfvxZ73WT8XcYzwa/3d7Q+ju5kLHYUScjnKpamf37Y4441xJcRYJNbBKNu4f
gYiuaQZ+tDh4WmOM3TDPdEGUpSsPAcIcXhncv1X2xZ4586RCEFMrGHpVrdTUS+8Wc/tvs7pDxgBN
zFT4UFPwicOmn2ICZWYio+oUoBhY64d/wlSU2fbFvvB4IPTeWlFrN6vEum3O0eN613fR+zHOf27Z
DcuNyn4oaTgQ580rPQPutiBWXNG+JvzDywdPrKnyFGT3b5dd6/Y2BOXEjV927MDk8Lx9HPyI306R
iZ3GPBMJbRxTCzfsgjW/9/nFkaMH2ZfZH6UrdbfFGnzNkFfIJVeqCVh0CslYkzENoB8ZT3dUt57M
uUmZwjn32BPkBL+9EKQINymiMCHUEJFw2tRcjeITxae7A3byLMtp9CkqGSW2/CqBPU/jVHN3wG2y
pgKSY8KlIkgBxhG/FwBgjJ8hxANwww0g473cEVq8GI3R14I2rbsABXAwYi3qkvHVW3pdeLh6CuPK
OumqbucX4j/iqamdi9o6v6PwyheiIwFVnY5z68DAnQvVUkZRlqz0NwxesiT8PwHuQrdpMY42dyH7
YhR27KZRKDmWi11f9xUPRqOY9i+lS6MFebTC6uIv3dEIS8AB1GAgF4naBtge6+2GsSuCBA5FOiBE
51uL4WVQUCP11I1InadKKjQMvUujlsyRygloPhF86YIc/Nlb7olhWmTXaUpPy5aoe9m7k7SehXy/
d8ycTLDhlW8Vug4QZNS0m1Venn7kZ+3yr7O1lMl4honOQL5aHjqenrJLJq+dsCsDRv8UE2Sz2KBr
MPun9ctGgcTlpDFazFSZVdVu4jtMuDOpkv/tW/cVVEOeRVNaxD1Z1iUQOomXofkK3+8sVBNqVxGX
ZBhsy3lboPiWauKbcRgLGVMcP2Lq6YATY0Is3KQ6qiq/rtGlhuKTOkmegB+XzYXegTCtwWqPjzr5
JBHW9IbcBvcwWUZjnvm3EipWVIGu39yDiE7LSsNWCO8vCeutPZPmKXGm2ED5YUVbc5tq+KhXq8tI
3TDQd/cD/FEfy/AqtaAsNvJgBYeYICC55XfgrcrUfCUjx8xdKuiUdrhGmGEIF3aJJxnAQuo/CXKR
WIG2ZmlqPBF1bwS2SdDf2ISkbg93NJKXs4pdgoKdINVia/FTA9m3xZb6LQlg2kIyX7cULNluFzbd
PapyPQH1PZak4ZlMQ4gTsw4RgYuX1Ra4E4dO5xVj57NFNXRkIzs4V/4h+cdzuToOlF/+ZN4kCHge
3uWsvEon9j9zI1IAZjB0xAKI9FtkbUZPZj5CXWdZBC3+lGLT00M1quB333IyWnEbE4ByGkrqK9KW
w/UUkvMir/PD23/v2ZTsgI+VOCN20UHz4nGauawGDuU6K3TgpDarCMR6B31DeewxnosEnWrrb0ei
3B7ulcAGbyOPE7yuuY87N2KHdw2Rxb9MV1CFAzQQJLTqgT6hRLZFxWiSYpRSSgK1BFa+F5g3l8Ir
tuj9MCWN6N10JqRFtolqycH3B7z5TrDM4TVNFRyw6V2cKQqDQ6qbbjHxYkh7MpT36pHXMwh7tgI/
WBOOI8j2/6/XYvA7HXv0RO3qvAJzDNEQpnniRtI2pyKePgGnuEq5U1MdjKJFx/pxaii0AHa1eOrE
7jGPKTBrH+5Tj7yLhMFOjltb118Ou3GDm+jYPnAtU340FMWCqumugDDb+QGMMcbW7Pyr2fNRQJw+
ox3jZpdkt+c5P9Z8dC7ZPOIA+90eQyR12uHK9UyCfqeQitK1Ag5fc73ZPy40mqQlZ0fKUHmDQNNi
Q8DpxasZsEheyxzkUCzbNtEseoDMoFquQB8Tp2tiKAyH56HtV4Okx3dahVOGMqCS+gl61f6cylAW
cgfypzaAoEqm44m8Ot6GnvrRtUlkceoAdRWIkJ3KuQgmAbPc9vJWeOKT0fjhfBQxG2ftW0/wOobW
132mrc/WM1NghP+se2Af8tbDYwFFZFaGAztwYCexy0LuGOlbJacw6vOpL6c5wo1CGgd/g2TuERHf
dVnFy+l4UIwfj1S56upYu7w01XyUuppHged9l7xXtQP0nE/lMvYPJr+GjaId5Oa8SCEYax+LiJcf
vN29B1GrzGRttbah2/T5itOG0NE5piEgUQ7oAj39V/65KMiiGktF4xLG1PgMhbhSaTESJh/zwSdy
JB24fQ1wMwRlRe940yFPpWrkH3zYU70WS3o9zjsUh+536nv36pkusqdB/Uf1Tz/zJ6kE/DuLMzOZ
RQsW8kSgZaFqKeyTBhk6xctZ6p8Z49cK16xB3TSwD0/7OhUn9kRWN9UZ7tQdbOLPZKzTs6k8GLcu
IbAdf0owrEwlIx8tOyyaop88UA+C6KRj12zW1HL972YAkGwFE8aHY3cB4ALhnIu6x1b8H+nkWRv1
B9G2QIP1StUH5q0YXgM2mpcGCOMQxjPmE9yetviBsUvWm77Wc8aQOdtm13Lz4nRIy5wbJVqo5ZsU
OL2Cd8ZGNSYUmjUX+wdGTjFNtzm3rFHbSiIz6yvExQLfeqlYRJZpI1IHCigOZT5iKpBVYKx3datP
55m3JFBSLOX9qFIotOpzUqU2id+7qQzcP3ZcQ3uJNdiXZH+68zJlqOM9AXoMZoLBkaot4374Jg3P
6ZhmVAN4p3ZwtCdplRHV4+lz9r5Gen5HsrCE+fMAEOWq1zelWkDYj8w7rH2IS0/4e9hWlXwxALxa
C7y0gqBcvt8XCCID+5F+B/7kRTfV+Wa4xeF32OA7hq+f1d4SFjs05GKx8hs5mtioLkW1mFNmTAGy
Gzg+kgo4yE6u4VrhESUk8ScNu3kFoqdHcwublVf8k/PRlmPFfrto6cP1nFqDjYAL99JRM5KLDyj+
oWZvVPrCWU5snHTh+ELZByhhv+7SvnxJSWEJU5nh3DchpbKk8ScOoazhn/BcYIZ1Sblojp6hlZjV
TMJjJsxzE3wK0YZKbTlpldpCPltl5n9vu/O2Q5tYpI6Rm37JQXVo504qqAm3+UuwtNY5yeqtXo/G
JfqYfXx6W1egwlJ23xYADIw1+1kl4sJ6dW+s5TXz7bdolAQnOMx3rVXIMNESPUpDpUOX0GPBwZKI
oN6iklRDo69+PXm29lND1f5yLLD2/5vy5H1qnSm7yZrCsk/CiPicjmb/EZEMl8dKeWsaM8KN4von
2Oyis0qW0JHLN0i83cYbFoXudvxfmcrIQuXxQSZTLM0ZPCPwRnkUWfXnDqjxN//tj/4DMJEh6yeC
uFb3BCeHdqaUuOadigkdokzQQBpWTqQI4WeSFQy6mKN9Q4l/MhmBRN2IwDE8Z92tizN1EePvs8vY
loiYBcYINdGtLzIiIGSwLWm67TKpEyIAEi1eIAkpAyrzzNVRN52WHbDYFdhLxFYX4c/UB2uqMKn2
0ZXfOFY6WefHKinHfTIevBu3Nhnby+ImA7tmcsYKlVc8tM35nuG8zaFjw+s8NVuxZ4uZF8epSab5
/qLg7cQZDZlMWpNECh1D3GzPdT8EFphqZQD7Gqn+ljeOQLim7D9qsEWJC6wR6s6ygyDsC17JNUhs
t827EbOMQEPeMbtvNaPlRPgwGkh+w+nrN3ht3dSCLV9U54yJhRVw7VkAOezco+w+ebhkMAqbQimL
G2jp0fqlNAm2VpiQr8dnNN7Ogot+ED2GQUptK4Y9uGZbER4YL2uFedBgpOoB92uLmB8ife3GTM9U
ugmTRQ/pbgx6jnznKTdjVzuNPllmwlcj+O2u9e6suP+MJG7aUQ7WLe5dk4Itwyog9V2vCBvYXAa5
uQMufyOr2DvqFTbBL4H9wu/t58lMu/kQ29thGCwcJyweN7JGS5CMac/w403ARBC1zUOhSMakg3Y5
qKLLE41XlZyUA7dyEsCvdwDNWaCXMyhtZxWaGMli5JDQ2SddXJ1zpknoZcPKAiLu/DaP8stWNn3Y
fC244MLV1GZtqTYdHDlFzzdeKszQeUMAiXfNpofmtngUPvE01nGCz4a8ImII1iGxNByeSHxOl/tp
z+ZoFGMqTS2NlKJKVmt4YOV2VcBOSrlt7SJSmGDh/hL2hOW1t1P5YeOqMxUUEI8fiwmVzntogyaD
2uWqP47Ae147sYSPbgO/kaHpNdZkq1e6lMDOkHbbChlE6xC85g65NwJT83Zt3aPe5B99cbKCQf/f
baFiOjNRvH0qVkHlbqt11BuzNkzRxX+ax/psTnR+PEWK/GtaMPyDPEkk+ohVM3iZeoTHNWHeQ/1C
dLMZUroZ5FkZ1SnCybLVhmg1cMTZTjWpC2Be6wB5n8Zn2JYlI6I1O8335UFVEG7JSjcOV+F2vstO
V5/iH0f+n5yDkw3mAjoeAvi7mMlVgYRFIAzYEjvWS/bHtMqS/AH5lTh1la5TI3UcbolVxPLBLBEz
nwoNaGw2MUfbCCEMPWAzFFvtgPFuirD/RqC6Rne2umxp3KV7qd4tpdqhy/k6o7XNutN+8QCQjzSA
JOM/12g3CoBH7MK962LgB+Q4B8p068TARg//psmr7N9eYli8CnvXQ/qJLyEY58FcfZswkD7QWRkD
qZOcxksFCeb2a0WRUVJWo1VC5ayqYojcreSpyOQd5CDI7y/J+UAxAiTat3T0uT3ubrUFc1lZlfh5
yuk8Dkyq+HIAcVDNPDRJ5o5C3ZTsSABeNzyPP8qV+vX94FdT63T8NdxN5zaJqeCjOeNes2ITEFuY
lmCA60TMM2ZGIJU/ASJ9z9pPt1kJN3urT55mvE0qAn3GK3yXyiIygFKzp2CDWzigCyTMfQxOOn9t
vin/+ZV9CVYEtOsQOcx4vGoK9k1IUArBQ7UiJlpjnmqyryIBrA/QkyRysZSEU0qTxcRzyKYm2ZZr
vLoCyfSILY2F6HbRORhVsIJLy9Pl4NyNofvyLxPWGm/hI8BAdAqQi42J5Q54ewc7zA8wQzPWULej
E2IjU0Zmr+Lc1xYEm95tf4g5xsxq72mEMeWzlBHjVQ29aGuKBKMAQ5tuevZRYBMihQbUTHCcZdzC
XuFBT6QEBHwKwtmhavCK5wO1VfXA14xSKSuU77H8fdq+73ZOWYP3Io6FONY6ixOqr2wTsPGakFI3
L2NTK4Kszlu62nLzsnXOHbyi+fBSup752heOxTQLXAiY4Fo41xtQHJUVEo3ai/Wd8Wc3RGHlPsz9
FeYHW5nbo2QY3cqsEjPEejonQy56pOJI9bo19RhaSA8oWAXfe5A7Eej+4nQ0WDGOHSv+cOTwQTBD
H249I0lUiVkCXrQbsV1F75Q13qH1AKDgIaodLTaVvL8xGx0cQGvIrc4x+jsqboStdjhbD7szQVhG
h/xqxSIa/xH/F+9KwguNMn6R/yuWsysA9i1+sD0xN1KWPkYHpxDb92tljmas0LpymvNUQedJ0dyo
TJMyD/VjJpVqV6nAs0zWoM0mOQol0GTgQAtTQQxwHBzxlyQe7dLbmMQLkgs9C5m7szkF+JLN2oQX
2yj8xsR8qzjqFU0NJ4WnI8urIqtk/34eQxzHImpiNzsXXR7+CYYNHFqlvIi8IQqfg0T80UGXR4Sb
Q1vSbmX7i4Y8zMKv6m6ByKd7ZTp0UGpW5+HXIVIHivYOHkY0cYIkfrHRDzMCHhO613GpNeT0p9Ld
EP1kpM3rvphsiAVvFTcy6+qB/QgqRdOqZbmy9oRnd4ZfzOIN14HGtLgdnSUVTU6Yx2E++5xXcs57
v71X5lhfjcVKxRK+v/eqCJAXqueNODKWJ+yfCPPrZRj/wRHchrlipF+e5lZ/3O2V9Utwr06V6064
VfD1A7xKZBk/M7ugRYZGOggdOH/t07liOAz4BOdQ3uM+F+xbGD8ts8uvDwZ0mh3NE8m9judySuIH
j0Fz9uNmpBfzYQOlQQFiPiY0bYRTy0N6DCFZbIZTpzdq15+f/4Rt51HMEWoTnONENfcbcPmodKTs
J3iYlmPa6jyHVG9t6V0G6TnHveNH6NvSyGP2XKyx5R0f+eZzi9mXLWH8V2DDjSaRik1UoLg8Jt4b
9IQ7WUfn1XMvxNhK0ViqDKpA3lC7YMC2w+HH4M/9KbggRfC8wbBLvK2nb9rWMOoKYUoJialdvL0F
//1hxVd2/xLbvQtqhL/RnOKRVGCeJS20WcH5MCgtQw8hFb8WzpsMnuEAdUmtoYG9cIWw03IpNhqB
HAW64QOVy/HICiSKG33qiC3LBT3ms9XQzTeTxaQYTa491eMnCxjycRBhgtt/nCmB51MnpXxsvuFk
SDWOsirrrahNTOLY3kjGhXvNZ6enekkGbdP0Tjy4cV3rMEkEq3lBbVRt3uUVDH2N5eLx8oMmxnwj
Xa+vnCtUtPg2oLPjO/HrCeXuF6iT0gEUhsYUKdUpxmkMpOmxqkRNgMW3nmUXBVRW4/L+1w4Lhs4r
RToICS5FzbWR9vbZbj63iJlhMEzMcjQJu4oRSTDrtbFCMWJXhz1esmMq6jfJQ1Dw89riiUT0jYBV
eCelbej1JACLMT4o8+4FhWkz5AjD+Ngx+L1Vun0au5JAFpyXb5iOJn4I+fsPOeIjZxdH7v3T/h3I
jokN2u+zsHo8k6CU0rxQnmzcQQ2fw+eOM6OkLzsGqFevwJiGyLg96scoSsst+LsV2uBmmQ9OTZMa
E99Uc5J0uckDAGr5+HBSlzETVKbRyAq7Vsogc5VA8ZiJp2S0X93+SpZ73ihSyrD0a4MfGom9T3N7
1DXXhNNR+77jK+UgLiKT7DVM32QeQmkQhO8H6jxn8JJz6rWZLXIvzcEomePourKnb4o3hWgfwChZ
wUp8t8JJCbYn5rpMIQim+SXReh4NkuHqzgVzSsmxy4IenkuaKuMLJEEU0NUlxDFjtjIj2MhGaFLH
+WlOXdqb12jlAxnNFyfK6Q9UQDGjEnhidwfExRel/1M7ybz+Qmcl1LXtJvfLD7XM9TgwmXVutYkK
VaO5UoLlr32epou3AS4chL2rr+0EmASM1YHUzDvlauJ1gpE1jpvfT7Fdew2ik5+mI9YJ5SwejtcV
y26yzw8GoIroz2s0bP977cTJs5m0njdWXFN67GHIaZWXIirfq2MYw5uMgktpIzVj8TLYruyMAXlm
snYosZs5TfL11UIJtoQl1ML+VPFyHYoKGj1TjrhkApi11VaTODnwd/oGHx5IlVLHSaDgVVy2ZOYz
FP6gzeA7EsONuIZCbBvdkmTcXpB/DtKpxwMQWvrxyodq0/l8JzB71ZT/3bVoDok00C+kPhhULc5f
/OSC36TjUE7tXTjaNxNvUgbWWqoUXcRxZRVOP2F0T97zLMzUJPFl8O2CqygNrq8W+TCh61kL0b6p
qQKq8EG8ViPVib4E2dRcOHVOLG0+SEsiTzqzj2poSaZtKVTPKizvc4cFyY43lUwZbEHxog0MhK97
otjmLpHeUuTDhduiU//o0OYMsCcqv8YceA3vW3zb+R4mPam1AeH6otiJ5I1rG+fyACsZfL5BJcF2
i2A1YnuT0TCkn5vmLRTiSgcfbncxpFtM80bZB1Sdyo2kXCTIIQy4FE2HBnAQNChSXtunobN4K+yV
9VI1K0XhGt9nyDYg8HtNKc6M5qROiV9Fgitr8naGtTS14wE9rQdKEjxFKGNYpwiTd0DzFGbdxfqY
UtDyXskJMU/7dSO8usPGEV5fvNvit+iKvPDD3wOj7KxEBuuCUk+AgdzCDfAaqp/WuftGIHEHLJCs
nHXrgxIkT4hkGRDLIsvgBloEde9MzK9q/G2a1xANNs2Bl0T0SKxL8K9ew6VV9OcilaOE1caT8OPu
tSd28i48GISCATdYVFZO56szfIbcwcCrDD1oQlvZHlvZnN7R5LO3/DCt9+X4uRkO4IN4+BbEVYeY
q8pWSd+A3ZX2F6QacPc3wezxtddaZg3umMSKP0Fh1SLS2kvPwONaI4hKEkMY58aHXqpHOKqUH7cS
Npf2gSqpSZPeK2bDQr+osRRx12bEn88lfshOCnQLqfUcKmXBjI+C3jU8Gf4BzsdhM4QSIsHJPhAK
GdQzIzRTtkFuBxu1a4hmaT/lkedHZLDKzyRPCvwVshxKKdLZQHU/XLR1XG2B5WVzLvTH8jPm8MQU
VkNKTn2jTk79Q5k/I6YoGFBGzS/WyfquTKh5UhhdI4Cxf7p0Z7619TcO/4wHPaq49LfXLhspZ93S
nTrCvuGJpp2BgorI9WuyLcygJdc3ayk9TOycCFBaZ2CwaBIo4ZNHR5l41H9nvGIlrZGmMoD6Pvbi
h6cvTmC5n5IlrB2D6TeMPvxiKgG126XfN/GttW5jzRoP5Ap+30HbQfGanzOy0TFz9KtQWz5EUv9O
2V23LuIRxQSNdZdNiAhSFAs7zZTZj+VFkolZmVTQUU8InmtW+vQeR19EEWr2JFk8z65HEkhWxYig
etSTXzcRI0E1QnlEXYM/3lwIGtNubJ/8G6xQiyL+eong7eiZdoKku/GnbphrNI77Djchwukc0pPm
Fvq0IcompaTrd7XwPn/ElL+Ob3mL4vH6ULXcFnmk9wvT0WZljGKVie4u285v2XqoGnUDAA2MktZG
NkrAkMG3F5AlV5hB84/nG1g4TgltHg1hoMBiwfYYDwMYYwdil5gGgYnRHbZgavamIJT/tCzwlnTA
yrwoqmhBnI6F1U90yXEbsYjN4ulGg2Q9UadJurehtZ2wBW+zULvTtr6bhGY8JHhk0BH/uhtkabBw
cEF+2ORjqjpVGaAz+Jlftwm0iX4qFjaSlGTNWbkI+l70NSDhgQtUF6aSXV1uB71r+iv5WgcE6MH9
CUChHw4KmfilFmPwLvalDQp7DE/i5V5HdQ0NgmASk+zLOOvVBBAJq8n5cvIkrX9om63/tFXjwYgl
TBuEJd+8k0E6ssSfbeJxhU5SzTLclCsWXXvU+mntQdBgcKkTo+udTBkXTxYSGs6bwQFW1tcE/baR
QcRtSdjz8I0TGDU/zA+Y9t/Q5hGKDNXIv0NjoGQKXnubldUKamnKzmg+nsJo7wrJ+5LDU75zvc4D
iCO5PJ6BYItN0MzU690a+oukP4uGlDQdgVYQj5zRAc5/Q6BKEvGe/osx/P1mi5NtDOcO0Aye9H8L
TG3aMqpPgxr38J2EiMQr6uv843wijoIgqXB6rsm+6z5dzwRTiJsjQ+q0u9V5tkQfyg4/rOZ4udSG
Dny5Cq9Y3hiVGcUnpiSkb4vJzMRmBeZpbqSv/EPdty/F+U+oanNNOZsFlTUGkh7YUYzW8pDYTTwK
41O6DuG+uMBgcnYtiP9bbrNbp4gFDw9u6PtoRbWO4tm5BLSmggoV/ArWXHTc9/vjbdEr+0LobmOS
kegJwpG8Pkud32WDpRqAhsK68I9QvQW7wQbMeY6H/KVhBxKaIxwMr6AKJNY/hgx2A9wudsPQqY23
hMjFgriGm6DViVq55UQZvPec9k3M/9xSecMllhVKwLvJiv02WoRacNJe5pFcwS9aH4jvkZAPF4B/
vgSbscF7ws1klTz8oHqNj2n36ZaBoMmggYEpNO840dti1A2FR44iz3uk/cMocI3X87DuAJzf9URU
FQqAuKfZfaZ7PyhwVcnum+mEnh07/em7WMeXr+ofaiccu0TWQlA56+SrzeFaVNbGU6KmntJmHay+
RSECnzYAbtM7mXNo0JJSPR71XJkE+yfeJvXFDua5oMJSfMaLhagac3acHCPYPyl1V30c1Znm8GhQ
4buxW5iNzV4ftfIlYHWVaCxXtBwaO8Sz+3WFdYK6ygYsLx9d3tuGyiQu1v2EZx4F3SxNy9UtkJT7
z/PBx/c0jSDgE6C0Mjf6yH1TiOcbogIYdPX2kt0hcdbT2wy0qa3+Kfs7YL/CHNeZKDdlFatpkdGU
ePl14IaEo/hoJuUhtnRSZQaErUXrZmLlaU8Xo9He7AJd5K5HqyMYKACjkFjeAP7lQbGJTbhWri/P
rj2+ZdFHpbvOUM6ATEQKGmKt6J2pfvl3XyCUZMPp0lpun/taVQe+tXRGP7OCBHTTaZIB5SKVNUPe
ME9WlUTEom5woUbT2nWw3FyNGHp+kF1UGoOoOwA/y4sSlLRCPt5RN4Txi9IiEf8LRuIzQnd+CLJQ
mbx9J0PqfmFO+SrW0KTNKv9MHIy0jKbYuLwYp3T8CW0h6tPlDMrexpWF8UywFbocZdweq8cYmY+0
6T67ISufwZwE/8hAOCPMu3SX1c6qtn36xErKQm6IaKE4HLuqJTXtfwIyOG9spas+IC0IRDhO6Fbp
d2vmMrzTYxl+2Biu8Ob3S+o7HjQB86KDb4XOaEeEjWI4+XksLbME1IRJSY9btQIgnKIwreJPjsdZ
mJ3I6ytoa+g2kfiaYq1TmGhOPLkksr6n15RlgB5G+W5kDP+TEW/brRo1obWciTgR6ixcf0NZjYzA
kkaWZXbhIZfCko+pcMRahWZi5GVHgsZrNdkwlrRaKxp1xjM3Vl8byoiCygbzStcslKXw82dYO7uS
3AdAeexpXdv8SYnBR8TXYQbpaZLspx6Iig6lj+H5J67QwHD3F6hgqA9cakDMvtTyhRw51NdkLn8R
Dh7uz+t2wzpbtx2wxHl+M5j0jWoynRR7nmw6GSrBWgV8id/IeqvobJmKY3HX+v+bqjRu+dFBru1R
+Rf56JEkNUa6YZWZy6O7lvngHKob7hxLrdw1vXjEmFUqZpt6zAZVLzeueNVZSgd7CloMlfDaizJU
jl/OODAJnpcpWZeb/woW3OWEE2eATLMXtM+zprRuFAvm+bhJ6gh6LtoC0sGDH6xemI4aB7E4Syej
j0+KT+ihZYO43xv03Re7ZwzZVQLb2RbC/Yy/pbOLHUcthS4dckdxQdSSZti9fyYKD67Bn0JszRB+
6TIhkrqS6ItzEqbZJ8aBvdIcTOYvF6kEPxYxIg1xEFiu0SEt7mzKmbAoSqMAVYf6o9T9wNfe9Yzs
J6LNqkCuDVqZUUXb1ef/GF3WVluvMQ2jPJs0JIuC1rLEmKR4/gaCDLeqfEzUklBA9afJlKkOWd5d
7fLbZBYLzhCjCYfB6h7kZpNEmi2R5MrgXUdU3G5g/CI5dUdaFkhIjCiBPpnpzNwWNa3NadTF8TW4
lWRQ+BzAs3vhRQRAfT2lVQRx8nZDmtRckR0mQ0PMFOJUOYc4iSxLZOAkE9yRgufKfhQ5MZr5FjWV
7owaKrMcQ83quJojiVCwDAQiv6DThoOAaHxu9X00P2280xV+TwDfx9J1/nhfw8NYxJqt4qeOa+cN
TvJ+Z0umBok5DZC6EdPw/KiJtsu21U9rEKeXXboGnqER7gY16bPQXw0+VcQ0DJ70noQiQLz+Ryxc
m+ktrtbfJDoQbGGhHlX3cfhC1/bLtBJpBDo270VQFGOlY5e9wE9pOMv+DNgyu8AYgOEPJV4+nnkD
Vh/ZAgbQS1F/W+uI0wZUzkt8gVdOXdm5+J/a0HGLufDysGekJIBYZUlV0D813H8O702gW/qEbPq6
lpiveVcKyn+Yt7RGXNj9qHAdG9610kSkMT/DYInysPS0VwWjrWV+5C3purKt2qxb48yL73c7dcly
OAic2FrfO81mlI+JDa69wYPyLxCm8jzjSOj9PIHSymHp4wnQwVxrDLcnPheTgiCW+7ywXiQfHLAt
MTUWcJGXeEbOsctw1jGqkJg9ojmc0JSeV6T4fRUm9SVf9DXx9dKqwGUNvPpw17p+gBjc3ZfvpV7N
fOQhICnOtYOBO47gJOrSr2a8dKqjIp+m9S/sfQ75I7Vu492Zt7+3w8DyBp0JE90gDstvVKieuaWU
zZgqsnYksKdU49/8i+3Ek+623u8YFR391h/oDtjqci3DC3rjcNTY85eW8KekPkG7eh3T59jKK9iI
UUEDJEBsDyLDpvPwScdwa+6ON4eiK0Y0Z/zcPaPMHF3GcPOG4GbN9L4u2V9aRWizkEvW2xOLjYC+
3Q+Ccl8HUzzidglyUeQIbnOukF/MJxqGG1CbfjAk/wgJRO13B+/iWxEdtk9awrfKI5y4lmBF9DRd
xVLUwaj1E4lIxT3PI+fvyR9hKR3AqIDGXI9xtXiRtojsPwmX9lAWRdmzy6xVhaea7lWNlu73JDD2
iXw0MYLd7AxGTq/E9jC8E54kHXFNUvaukYqw39m0nsCDIZh3RsUrMCcsFcXXBr4x/NdB24qVyxT7
tDTSVW6uIlGFcxfc8z0Ez377h1fPx90v5h3t+kWmdFjaAZE8n2uO/M79WCuMfMK/F7UfSiAtvo5Q
IeWRYru6p69YCLEcWT7ij72DNf/mg/y6gih2aggZQNtpVqeVUumAEYrmV5QJZg5/3hOh7ExwAQMu
EACFYpIgaCXCocs+oVxlh3YkF++05brcDwQnPaJOwww+nf16gvnpctK2pKUIs2K3toXjuOVgwmIl
2KbK4hKoNThQmt1INM7afH4TzjUmN8wQGQ/jmbozQVK3irsa+74lX5F/A5B2zru3dGuNV/NQAQ/V
430epJULwitzsEbDUSWVTaYZVbnv7Jfp7vpuRmVLVCuIoRzxvCfnZ3++l5IsvUJ5vuvRbtEUCmiN
IQLCdx/D4G25DlU40hWQtXftGkC89mgVuTQFpxwrW6cAkVNesmmuSp1aMWXrxwAIpsjWoK0AVwpt
wyI3yPxBpmjBR77wyBkK6EYC4GCrbE4nKi0k1nNO2kx7zNwQqOI0fz3jcURPqvvfuzUM4Z0skF69
FkIUdR4eJkPgYc5zuvFsvo0/bjHjD/n6satyDHKELYTyYawpuWJA7IXMAOamFxiz2b5Qny7BEN5o
3Hj3NmzOjoguj+wnq1te9vvPc5Y4LcWzaxSY7LG8lHwS3IMrCen2v0LQSBMqZoGpmyVcfMEbeykQ
VCik+KqP20p31sS3+wxNivkz68M/F4teqvK0kh76YP4FYpKEJ7fakRzjTdR7V/AukqH6zVteqAiv
fILsHaH2n0d5aZOs0XMAZLZsjhBJzr1L7ykeB+j6+n+slTf/rbWjS4Ip04StqxvHJYPot0TUTab6
GHpngGuS1gbu7vHmPtKgiHZXZGsUKpuGhGHocLGpNHDq55ElbBUpTmnYuMuAnN5j8sUAXo/IW+Y5
/W1v06AtQZkruasUZlIS5bBaVap9ybsC8IEB+JGgSXp58cSEvVboov+VrR2EPh4sd2lClHbzptKC
8em7jz/iAQkAUEp0B9iN870tghDeqc7vQNw2w21aKZWxNFhry+CgqaY8MyMmchMc7gmU0HNpURVZ
vbcP62WrSRX2qJ9CCYg7XSUB/a5w/p/ybj8e4OyTr1ULdTZzzQXs+MijWVbioVakD6TFfsfJVsGt
Cer070cM9DrKS7xtrjyT1pZ6fbudkPJNj74/hKOPfefADdnm91rUGv/tfBolie4C6e1ed3lnGhb/
psfX/MGIlBpfAo0IP/+lb04/8MpP6vSCakEVCPe4w0n0cJp/7EEN48v56m2AkEX/smAG2KQAglM3
Ahu1FbCArQUBbC++2AUi/IqsgG9dMQnQWajs7P6j0GuzSNy6haY2nSdUMUwHPdv5bHHwpVZCullf
TlO5HJzP685BelBotWXX/hBScnDqxlmtmHrLeDOVQPyOmIXva5trJBc6FDi7UpZ4BpnqnduReJf3
ftv3e+UZ//RhPCmwQ/Zs2QACbts81kfQox3JSwU+SE0YpWMgVPO8JZg9jQtAXGswINVLgND8Zb+4
iZuvonNUALaZkJMmNYeY3kH9oaNo76V1Bj+kf3Hl+21Qg5gwMj6R4mTPjBpaHpWA431PpBwTmpSe
/VsNLKGdqTrBXEVQwtOsPL1oP6kb2J2gOsbcG/3jGPwlw9zCHqOyd64rKkKcSPG6khHPRSZQdXQG
m3fK87f38qtkELRhfT/mxT/oQ69Pf9MN8hpqjNcT9wDNT0YULM92YdicQGB4PhHK4td26P0fLwHy
SsSdMwFeqM07Z/MhIf+bhcCJu/xGvLQmBifzUtqFNn2z2LE4Fy6MsrgNpytQma2uMgjBdvCmQ0co
/fumqdM/+3znm0Wo+2jQoMntf3mvdlnCC7XdbHOYZ0ycSHtaYa0232vvRYmcDL8FqVA7uqylaeYJ
MZI4pWFa0MxNiEQE8AQBHoJ+8XF9QVoChcSBmi1yHB1+2GCbnu0XOaNiXirwCfwRvsfLMpCgTZjF
lEFBCBcLW2ttZKMTmEUncFtr6nUe/x1ii+sL/2TsqH6J0f4SFbif34yJap/phjlrwH9pHd0SXwHl
dU2/qM7lCeeACEfdjr95OSa+FNhwPygKxbEHveQhWcN3aJpL0Fy8WEV3kVds1x24n9rua5DoLLwE
mDYT2u+Yvts0lvStm1LvH2FFvNMaqnBTEj2rn26lHnQjMVp3GN3bK3EEKNgiWHUTzK+EvLhARaoc
BJCXk8dGsdWUgzAk59Lp3pemwrqcfgL/0hDqik0Pj1jZIDhC1RQDkpO0kXAAulpe6asBlY5EuF7x
bboSyq4/RIXe7t/X5HxHCZQ4X8+0fh2oI+WMpTcrRJ9KhiqTI8ZCQYAIYOeWvnrL7TGIM30PX6EX
5rdFyl9vY0IJ9RaJ35l+5PcSU/rrE91ARHxNgPNn4cE9buZ7bHBcBXvYJCYmNdxvgvbf5JTPHsyW
eoDUpvwGPT0JoiszOd7W/zY9H8ZuwrQyWp360Wa2+Sgw2iXUyckfypO9w+kONHWGhTGyeAB7apGW
4R08w8lVAJ29dRKiS5IzJShrRkndCXH9rmKB4osY9FBbBM6gwEB8mWdVubm3WlpyTZnPVTPg2v9I
F5lbqluFtdCOcmE9kfVTvBtdGwuGuUg4xlYRzT9zTdlde6VtJmGSLP9bGWUE0J2UagvAdbmLi2vX
fiHTJmsLpvmwh3cwTcPgkdmXx5HGa9grX+rmAMDpoI+rNxRwJgBNzm7WQ5N0IUEvQ1nT2BSEcdv6
RQ6hLdxSVolcYmniNLAXczAltmd1cITzd7Rd4FhNEHGZNwyV90WVH6q4s2bV5afhI4RcRKMVa3SO
+Nsvf9M2RMKlGx1JZS4uZpZfLOdQ5tThf1d1cFejsDogcmDUacO9FWqNVHrJRZl5zp50I8f0Qs/l
ZaUQroKZsMTpbYQP2n5LXOjO3gWQsblt5Lei/Z5gpbrbBMJLHpzoGQRzEWoR9kEaQIdAcZkBtlo+
jDxU3AnprvmnJ9PQ6KM0/qmWdy2Qv1ibtJOF2/hwTpW8GoZIT2k4XMF/z8ayVhlPGcPs5bEpzI8f
pnKbNP3pI46JucdGZtAPUX+MW00/hc2yu/wNLcC4jfb3SISO1MHhovZCkYVUgVbIpWfRK6r9kGAC
gqgORNuqBk+y3VpqjDCRK9H0ek3TkdArxiX7+OBqWWjWYiES7SE0UTQNAS8XgXITL3ePGQ03fpXd
3AJjBkW4LnBUwEe6c0bFKT2xN8SOqaDzKBtyLQbkYPgolC9xwisBM1txGcVqAintTybYJ2lca63R
/JIJJ6yxj2jqiaIeMiwmXyCLN9GCScbr09PJw0c4bFpBntnsp+3yE4w+aeFWl14lAA7l+RC88r82
qSk3eqyUIoU+9f3gt7Pst01vLWRNBXd0SsV4n5z/4VERCbLvKgwgUxWFmwC1CSwNkq5tL07dVkZE
YQVNSrJNv01FRT1dWVkmdmkONJ44Dj0TgIujwV8MDzCZk2PQ34pc2/WntRvokvdkJ5eus5StbQhu
AOOOFBCyelUsFEEgVpF65eFtiHdbn2GWCCXTQPt7zXPUzxQfAEpd3eautfhTrJgw6scFe2A+kVU9
ycX5gHmVZg5XI7nH8aO1BYWsuWiyKmTsFq1JNR8I3quVANkOOpR5Jzc12dHn3BHPwIDnc9JvoWsV
72yIfuULRYftNTqHUbuROQo5oBSQktjlg3yPdGCrn9DkDhvAZzbB7Fdt26zNIg61eLzQkEuWPo7z
k4dyx85rtV7U2noLXG76um1w6crZbZOz2Q1EHrq6EpYDc0okYfMVbx+GucgmuylIcTlDlhbep9bG
lckgIfZxHsMLIoygsYC9xDzrxl4lTzDIwdr/5KeJtjpgyqZYEGucNyFzslcmSZahdPIXKKOoklRo
Ht/Ap+Nsz1xA+2DYaPWYnPiyWc1bzu62Lwg3dbV1dzG2im9+/ujH0Cr5gae8r6V+x8w42mFc4qs3
WUc1FGswXOUGcMDYL8ZpScxORLEIIL6iuBQyfpiHzP5vPSu4nsBVm5jJU2Cj6NAM1mnV9KMg1cB3
vbYI81CPzC4wZvwxl3iKaOnUZPYNphgAB4/YmFZ4/s6WD/0a78LdqAtEG0IMjvgSJ191ufnrLd5f
ntkpwj2JFCJPun9C25ZQ9L49R1KQ53R1O1n+0VEQc+O+7XoRWnjnvVi9/yQFS0dMcMilOMxc0K+f
3fOUYQi3diMG/fR1CvYXUmU5wEliHExRnMBWeIEorWR0O02RC5+mSVfEbaWwDcv8SotO/jTKnu8l
HclEPhSlw8JtAJRDMqlnH+Z5aUPLF9iaCwct53I9tvXScZITvm5CzwA+8M2/pWyFTDOZaFZLrgpG
VBX5FeDTt/7N8xBL4PukZybMPJboqBP4rMDDhciDc1vLBmW1yHz0PJRL9Vw92zkK9UPNd2F3dKfS
0pHzAgi2acBQ6mA0SFyp96BS7wjYro7sIa7hRcaCYVsQM9cvnDjA6umNQ2tyTjpejt3sTepGsWqN
148bfgDsPB7r0F8zjx0o91yCE81944Du8hXEN6Kaqf8xFRovWOp+ku7xwJkj0dgkAt4mGs4Q9VFX
MpiMZAmb5hWjtqYUDAEQVRwMGqIQCHLJxuvNWTv1Dp/msw5RZ0atAMLhrq41AqJdZGWpefRBBxH8
2FGmcDENwX+x7C+ZkQQbwZ0evFLupLMcsdqNaFq4NpfSwM83a6Go+3tQnCU4PtbvcPCrttIALhTX
ntkCM7WWCJwyDC1OXAWhJbxhIGK5SpA5GwKDziEgdZeurcaee39vegV2CyRqm0wmLcxRh+cXIgMy
ctNdiJu4cM3ZLNnTOFNL5A22AvTekb7z3P++ydREMp5vtIb6CAfn/CsPrMPCtzT4L9299tUJjuYt
BpoA4dlRdN3bdXCInM5uhIB8nyv4eApLpHieIOUYTJ/RamHtrkmzlf5yydZvoeEMOLIXNwvhGFgl
k1JqWxsIJ2nuoMoJtrSyTu/Nc9k1CWQsw5eupf22iO5uMP/lA4Y+esQQgCdMEVS9ekeP5jE67jV/
khE7WM5o0Keb4vYJ/sn6lSo0w07hM18DoPuH91rvbmQ8fC4Eq3f6CRCjnwCvFHZ5PQI2L7vLNkY/
Yz/2finVTHQ1Rjd1psUt51DpszXd2VFssk/l17x8FF2OrIbttoeC27GB+xtR0lXFDMoGYmxU0SpT
lUKx7apSte0/1pzC3gy68u/bPUn+9XRszRNeTaxZfpMdfpbowIqsUp0ZOTumMPKYDoY5JZ9CU5y6
EvDNdDK6nKBE6typqXoZr/SfVrZx15cdHzoJZ+GNbByidXPOfx/6YCBlal2ZMZtCfWLrr7SIOVjd
gl8HKG/kN9Vb5LP5s/9PjtFUUWzNfEdUSunixXlrMpq8eK9H6jsWVqToznR3aPbicLnBU5mBtN18
gjKOl4iw4FoCUiDIJr2HFT1hlpe28OOVPUYq3xZgoLagB4Ew7SR0Uc/7XcpfCBqHtXB286C66BTU
M7V+E81VO8UGmB8Duyyri1v4tiws75loRIyZPd+iIzpfTcrfENPj9ALY/sNx9GlNhFCc0/CEJAXO
OA5rbQY1LR/o2Y81kuy+MbZ3SxIs0aTXhN7C62XMp2875GKDzFOtVXjRXG4chZ5xRrR+Bko1ccdX
+tZL2DMBRKVdIUCuaybsLQRUJr+ZKToCaAlZhXPs6I/RcANW+d9x87fANBBOsR8oWrp32VHSnEiZ
rKpZTFXcQXy6k8m1TTtf8CPUzIFtLakrEQ9Lk6tZytQk88RphgeFJnjdAuUFBQw7Z5QwXpLkqKa5
Z3rf6VVgtoka5Wdo99Di3x0vUCdB2sfYrrYp/1ev8h3agCdzdsCSj8qmLDLOCqSrIdFb0Y4d2GbG
THvEOzzgNQ5ky5EYsynSQ47AfhjezVd5ou6+N2Fufeq7R0RAOjudv/GekNX3dVTXTl5u9SoGdZJu
MlxNbrzI2CgeCYzHznZjlJ5eup7uwgWvarkbsGRMbdglF+cG4Mp28SOKG9A5DsFVmexm9JQurbRr
xZ9jV/qZ4LPDJEjUGHPNB28WFAahI7ezscThNwaj2SfQEClnB7tXKQpAyg8QZw6mm3DXlaqAdH37
7FfuNyEu9Fgp3skKaY1GjWAA7VrepfRdKFx0fqw0tbzaJA9GX5POjcJmzU1Hm4rpahI/qNvT5DOj
vjrhgUphzqnPQTm6fsdFZi4P7gCRhR5uma3/MRzoUpIv4My9XeaUlLsPUtxR55TIprO5yEF2t1/1
NVmOhyXYhkhA77RRpSuMHcgHXPc9ekPh+16E5gsSbDfdHG4AmdCfDMd2ah8jt8/Cg6oDOgURpCju
VBaq3Kn71n1fH5rysDZvnGtpMXURc31F/y2rE3x3iJ06oAtXzVMd49qBiOw1xsaSeMQJjWpCqUaM
BBf9AXWHKvpmSQLXbERgmnt15kYy5ASZdbw7mMn6ikz+tRlPERq9IOvXfaXMidGF6c1YeNMFFW02
CM5XUnSQjJH/Dsv0qL80pbF1qDIdhLqAVNAS8xsiME3z7go60HpQQNEsQQ6g7Wz3q/zeV4Zhp6ko
PJBy6FpK/UgOBvZlsvG6+RqDdEAUoZMej1bQVR4srHWuwm9gnhQp0T4G1B85NonS2NW4gtySNKIt
m/PxZv/09QS4ARnfmeiIiqEOEcy9VxRlQKrDXLVAoZK1/Ldfnh3wRzI2wsmZwxWGloLKmphjJfDM
e9pcSxpvtzXwGmoWU651IfX434IoUty4w7VZOnMC9y74vDzDVz2J+uhF3lQQJz33y3Ixb+ECFBnI
FmnvhsjtH9WLziaiRIymfgvT5bSuFkN5SxcfclxviXg5t1ML+vqku5Nf9fZjdf/LfOPOZ/RS1dtD
nUiX/aMo5DlVeTsdFL4VIOM1GF/SddM1/kVViXXEPEsyD/wk5IaDQzx5ENDKORZ3hoY0hFfGRnpi
ROazjaxMRse2dZJW9ee7ydXRQmvqB1JTkJpBLnp5TJTyqNshurwBNKXXq+UNj6qNWxArf5JL3hUo
FQ2YPc5KLbLpyIXh6CWp8w8w4ORKk2Z4wm2O4w36Xj5P5JwRLjO9uXVUzmSGjgYenaJtTt9B6Syl
jjfaeBqmP8b7sBcwL9fgA/fZ+71tjsbxHZfzfDccBRqiG61fdAOP4TCI1DZlI7HnVSFhmsqgXiO5
Jw7cXfFSdXSWOH1zfAQ3n0/B2DsfoGE9+FYLejp5qOvhp64n4MNOuDJQMi655LuB/af2ZErZyIZO
OhfazEdUgH8d1zxMbbBPwW38otnVfOjjO5YZzZ1QGVBxAnEXuQOPwYFd4EIZJXAm8R1R65PSys6V
S09hARel1NLqQl4LJCcByhwrSdyWiSzfNUaNCMie2xxGdrVeUAyXBbvdWwn5LpTFqGhXZwJCjmrv
A9o0Mioos+2rWk6QnPmpFZvhFrKmNwHP8lZPzWjBz1fyFl0S5EuSHsYAOM7RL4tbS7jZSj16J78s
k9aP8e3zM4T+mBdNbz6dFhq07AxKPtLznotaFqkbb3NOsBFT/TxHnKMrWCqyk0Qq1YgWvDwumRuP
iE8dWcXJtp/IHd7VXBwtqyXJGgT+frfSlKWSk1oZMuswWDc4TZbV7KX9rVKbPJsHeA0lbWAtqcmx
7RuFChqfAzr31ds9TjgRNChzNJYQlmr9gyG6kdVPYbBr3dW9fBZpc+61yh9A9EeV5CQAGfIHhLbR
AILrlHXfvRJkRuyUxM6YfpqaREPmyOXSu6l60zhd2CFW11BYo1W3qiC592fNYWhDvzNyCd82PFKc
+dRMk2kJZ+IYMidDrM0MxerOPT/1AukO6vMu6uVsSdQ4LQOxML9t75my0jKCzc9OOgTpCbFCBWR+
iTzt/t2WIbkhcPTBRV9bEMLGCtUI6M20WFoHE8YK5Mfq12fhp9SrA7vbhKmDAJhUGVpW+jS43NMI
YeJae1zXaWLMUM4FIuXFYFePaUjXHFMRZeQ7Jr86/6o4d8B4pVBP7HS9UkVXc09LaEVT/Xtm/T2C
rH+XcXiLru44laprwZVA2XXa382K5xgT19Wwx/Qyw2Ba8bVBi5AaoCxFgKTCVbhhxDKQoSeeHxA5
kuEJTCJ7Ca/SO+NAQ8GHt3htd6UsN1ELX6KQkD1kKGIR1iEC+VIYp0PO5jYgDzunMxdOsVtex6Wo
hpqG2AUBh8oDsD1eE06d9yMk20/edqF/CIkWKLfHthq6c/nWwXKDjFJdgXVDOq4vBYf0Mtynewtb
bLnBGW22Rysv1Uzw88/SY2go9BvqakdDQeqSjAkaVifOD8VP/l8+Gpqvl/9QUNGdSd80Z460A2Gr
SjjtoHe1HZmFkPBEpxJZVWYoVnFIMm0Cpv4sB/kvrIk8huHeO9b/+2OLci7EgHj2OzEOokxpeA6d
uhMLz3mLXKux4raY5RaxjFlmlrjG8j6GLD9wVQAxBwjXcXVIlyeOrXSTsikqEU9Z7oMIEMXXjssH
l1LLaeKeYYKYzlCuCuTlcqeemadAY9q+mVNoDjWZSbE7ADNSnXlHbsP0tPweOgseAVExMniAfNiM
RkYqRLjGMDzC0r1WeFL9/DEdPxWO4KlzoLwHXBnIWt7yp4BpRGXgIbaLr+5YPk4XLUJ2beTkrXt4
ojMLnAW41knnKMIQxXU5PHaeDXZUUU7zsAe/Tkgt1kwl7cKm2R//QSRUGfOx7YeTc+VWq69hqcFZ
F+mi1BsDnu17uZ+wbgF/D0dVL7t6r8X5T56S4ioLJKCIMDi/hmuNHWxRQox3E3zNmOJBZ/rh0O7E
VvYagz1aSp8n9uIwUizqQZYFKd4J90Om/W1rqn4MvoVJdg5dmrxT5a4FlQU75SmCmc6c3pjP8wN0
7OOz0eIVL0jqlsumViomK/DOjxzTI3TW7EBmSLU/BZ+4ELJ4jr+2F+c8xviRrfavc6aLMjUS9kTz
VZTe64gitmhuJ8j2BGXio5l3K1ztR2YTt0eiwDPl44Y=
`pragma protect end_protected
