// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:52 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hPTtv5eJAEez3uvlkH5/poV5hrPf6wNhJCW2nt2bDsq+KoJm2b2U8fSprzq3+4mR
4yIOHxT5hPVIhjkR0Y7v9AQu26yIHdvnL/kLbiP+GP6uptcjD1XGgZdgRvr1KjZC
JNAcOBcWazwZXFweD4W6Wqnx6xKpMALroUw/3IS8hro=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5568)
syll38vGemdkbpv5DORgkjlZ9PxmiqQ+k2LokL6HkMZN5uKvseIRS1kWAELAU9CK
pGkPYXRXBXelGCUcwRkug+IL29bp47avY1f7zpAiBwkXQos+39mvIKsytr1OeTdY
uFL4IYD/131YZL39hY8X3Z6sgCPAzOpW9DbjvEwlB204qMSCd+ef11gBDYyc3i6j
d/lER2kAj3YXofeJy0auqSZOdgHfxUV0w9M3AcYgtJHFXR36VLPZl/J91HjUP2Ep
Qx3ziP43zs/W6LEM01SZAbkgw9ZThhQIA8mmS34E71G34bC45f64s57YmZdtKBl6
RW3oV8GNXEtbVk/ig0XZEwqWUi0xHsaUuKDu6kr1Q5Xp76ThcQgAt+kRNqYB2KIu
imbVPV2vcPba36eO7U7yq3HKRXqpSMLfjwk93LneIXpSJhb1ZmRGIxDsSFkzk3nH
gjTwZGo67KXykkgnUBa/BFH8+l0W7ziyw9DzK56X3kezqhMI+GpIZo8boWYHt2tH
houu1X79QOYUIbqNCYXxC4pP/GeuRDmoQ3XR+OHo8Uvi/UErBuzoDeG0wspuOXr3
/ppqdCEE+dP8MGD0khUXo5HmOCsqwlzCvKnWtY3kREFcM8FU56wecR4rnHd/bYke
WT16pBbuKDWvH5F8KsfiMBDDiZP1jnvenNv9i36+9kMEf3X+bTeeN2tO3rFnEPVt
cnzbA9QTCp5yXf59nAxsxIO4wZJE/NZqXYEjTwxXS4bHzy1NtQj2FEh6rd6/onSj
EEUlvDPWah2hBKq/nVgMelMojbFdBdyNZr0JFBCQPsaHlaeMXWqFTQbGTGgpqeLQ
AhiM3sN9LuSX5/pt7rV9hVtbHwBoxgT4nlt3prg7EhOmAjnd781h5Ch0tNyOUYUy
gB6w5OX311ImEGmn4UtVd68aAdS1eGdoDJEVKisWrUDOQeB6KbnovW6lVH6oeCCE
nBvd5rseLzrolwfXrCUBei7fPy+WHx3QQuLilR/cTXmtiHjEr2aj6E8meev+jkNX
Wobp/p9s2ai65+EKuNy+gIGRFsglrZZo2wKKua9MSwVnkr34PVcJenUTH9uOiLjk
KFbPKRAWm4eDdjJedoGktQj/A1EnW7ij3ZFFI6WCryERm0ZTUCahsQm069CikcNP
KULv2Gxmgbj7h3QBFrP/dLAZ0oAEfDrbiwCFrKOVmS9j9lFwQeKsAMWncWLPwYe2
ocF8B0edOqbHjlbgHI+RQ8ay4E3R6FZVZqu9FQFvJJXWI2TjO3VfJgVSd3bBvFMY
VbMRLxDvUVqUDQ/LoEt0KeX5KhY4b5otwM3/1IWxa3eCTmxcxSEaXUKyWQMrZR7q
q4lv1MOwiGfckFB1VhfgEf+4vsI08T3CJUpFErOcF9qGLETAU7tSold47CAATF+u
VHwRVWR/AR+sO586nPyHNl64zuN1Xbc8G4zbHK0NduHWoBn9PNGVRh0I1LMmZVgd
ai/dUT5UkiANzVnP+4BzJ8x8yVF0uSV7ugHVclGFzl2O53LlcmRc9DYxuXVZ2g7m
ARD9Cmq2ITO3rR0xHtJl+r6O6ttKP99egIkS6WqZnlJHxpFtc7ATcVc6HThVO0Tv
ZHJYKQknRYJNmsJFxb1oLXbM2Yg1wY7u6d3O2QyGF1JMfMoSbTIuUiBTmlkQbRAo
aReizCzlvhsfIWvP5uMD+i4k72DdKcgEgLMx5QzyezWw6SbEy8iviEMeZFt5lo6j
HXW/f1KAuqQhaxoZhFLLiyzzFs1LkH8m+RuCOGUR/R8kxkY+5Oc1Np48sx5vF1lJ
uQiDhGGdr6MHpn+dVIuYNjZXQV00cZxNBXD6MBJ6mtilSqgBIZh8hLSdh+5UsbSB
NlMqKmpOLYwh6mQQK3VavEEq/b7c+/XofO4jK6JMbQXCELmHhz24k4tSZu83+SVB
T8IMC923/pYVexnTCjLAjRqwWolqdRy1yvKg2cIOiJroq0v/LfqaAGWoLmfWQh9A
1T1XjcD9E2oofrXIxRTel2cnnHL3cTuC7NCyN5+H5jhW7chFB1DShGwAfU+l9x7U
dDPeykdH+6iYBMCKJwmd1w8w1TU69F/hCyLZlku7d+E9lxcsjTkT7B/UQHC3g6Z7
0VbdK+Hxz8iYg3S2ShDFEDcBa+OlObQEvAaIdjrkI6Mv11Vu4+Gk98gh/HTxxmvf
S+627eFSl0U1SIJnodiAJHSzDEERy4MnVwU0RTfsuu4/TGxk2j21qdmVOS1hBtGz
2sEqWOUo5FlEY1Mn63S4ltkyTVSSnSZDp8beHmCL0CkipC3wt3X7xp2zZAT4/hnV
CQb/WCHnUJ4/pBde5uOzDEQgZjK6l1Qd/c1BYq76JaxkQxpwBSqqdKLIH9XuSR9+
/O5oX66bbzF5FDhtPkOBUzfJwSano2pMp/SeJtpS9kmlRtWuvMBVp8ocfFANEwm6
+gwvs/igKeCX5HnXXOYWgYHBQowh3a6IonYiL/YAqUt55lj4e4Sb2gg/MxOomnYc
nTMJUx4CKCrDwtsiN3/fo37Rxx+6MqoQNW2wWboTNpi8JzfxVe2yW8agkopSNiNw
bhRKnGV+Min2uxCopK7S9dBISBX7nwkna3KGh24+QAgBfNIUXPP6qz6z6hakLZEN
6Ao1IKU3JBk/4bMYPbZ03bRhu79P6BagMeL2sezD9aVLMRvopricCULHYRHESBL4
UrZTGV9lUufnkRRnu1QCTUh4YLB8/EG8yCziWLubUKeya5TYHxp2UXWN1qNO6kaZ
RrcCeklyL+LJfLDvcJEHrtfcCvk3RnaINCnRT5+jZ6mcXALGb5vzdHqtb0uNdCdH
H/aT5uqOkcf9r7FaKgfiQafFaAp5a9c7x7gjCsq2bu0hN2VkAfMTQyz5FxD012mh
8AGY57CfYLhL/5gqpqhD42MYhvii0fG4Zg+LXRmC8mf+udn5pLeS0R9TwqGuTRuh
jeb0kfb3w26fWSBUMcCJuCOBr+uL28eekToZ0M1Vn/lR9b0xT1DFrtkTJLP0D/Gg
zDzOQYGANzu/Mavs63Md14jpscB+dIzvYWz/r6nEiliu4AvRWJFCKg8bY3kdLAOi
H3uxXSbbZKcLi+Ne0Pkvh3VGIJ+FuDvntm0ACUOjUJgyJAwQsz0Flh6oIFoz/CB4
iNKNyZl9/VNcpRcCZkqEzbFhC8BgTmJB+F2HPmiIQrE7xeNovJWSS6YHsTo2++s5
0OxF/Z/QHXneo34zCblIlSKOVsewPfVVbgjivGtTxu40WybMWam/tSBolC4MlgGQ
PM/3iIdpIWCpSkcymBRLAKiSV7ctoEtMw8ZJhIitNCdG1jiRbVI/R0HmCxKAPOec
LxC/xbE+oxaUELSgBmA9G2+wyTZE/I2L4K6OyVsKyZR8khWWVQ1QGudsRH9+fASe
2mXI+EKLp1QeuQzdpxZGml7SR7E9feBhlfFrm3RkSAuDu4LWlgVs/JkUnE2xXdSa
rJSVVf8+CtdBaM/YH1bid5Dj5zdmtXE7Fpx/cUehRLR2XjySGxwMP9VA2skqqGzC
u+eAEgZsS1W4OgrZuXPKmmCCKJe63WLYvtL6veC+/fksLG3smcELADpUbBr8k66n
FAbtPIllz2CpMdE8tMjEYUYk/vnDJ/HCfddpE9eQPKR/ZLRsWJrrQNfLojPM4yK7
KRuxODnvbv032R5GbLScHOl21O/WP7C6n4cL0eOT30p8AcKcxIVIbxhUgm8PVmLG
Aj2R3fi3BELKP/1BZEK0+LXKlDK2WKTGqmqIogYHeG40y40Zr3BLAdymoNP44YNJ
0egwnRWvpzgJlcOIoZZU5B4Yn7Z9xdDazUbXJ5u7UVpLXOL0Y8uXoH1ZCUlRTuhq
pTUz/3AUjnKTloKkWJ/AD/NIRPcTkREOV8guNSR7otro7D3o/p1TyRiSwL98XjMM
Py0+6VCXH38F/IzWqWggpsDuT9ZaU5+ttm+9vUwj7ufcInrIM0hmYMCV0hTrjvIB
uqzJsyiddJNHpvvRW24XAr+6QaZC2RZpLjo0TgU7n3qDAveWyZWEB9Znxd17j3E0
XCQ7wciLOdHLUkSj3TPwHPqfYcjZT2fKJpS9wPaYVcGRtsp8XCyKPVhPdkJPV/ve
T9IqHKTS9236sBIN9726I0jb/YhR7EYhAvgh6yner9RAtu/UGryAB72CK5D6Bhe1
0CycHa2WeACxQfKeyaIHMQcKWCkBKvvYDyW3SfwV28XhDku0B9UFkLor5V3EoZdT
PPzZGIfbfCG7+CjEc4iyvElquZQvDF3x01uvRsf/Q1MRKN2Z5lTWWx3+q3HuapMv
4TwKxFbXLDxomU9T8B8BDbPF3OtU7xDAhRfHkHjrz+FMNcROGVZSMhw5dAP0mL7q
AMG/uA9qwkRnmJK5P2hyjsJWU6nPfUlTKKCXLL+sYDp1imPT3h8/gIHIrdcjxtJV
fU5Av7M8gswby08oUi38iz5cxMpLd30laKNEXwEcrun6oNl7yKDye1fzq26SY0Fk
UCp5iNp9ef0w6NFPqZEQEe524LO4M6voCwDY+JMc/J5mVZRfGxdLX8+vexBVmZm/
INWpQcYrT/dp/PVYVHvc6N0ABXAkT7nNqAAvN/aJlu5JHXsHISJ4gBd5cVv59QJM
TLMzjCp4ODd1KCheWYGkjtNJ5ZmG94wFFpMamGZkTTjX9pDrGhyxeGENcfQsS89Z
GTusXjP24ghqPbmSn54XLJQoQ5f/9rHxQFxv6uyAwzk1nA2GaA8peucRLxfkAAKG
JW4ABq5wWTXSH2zetRgN549pM8+J6JI2VD3KNueEjwMGN4Kc7yLryDltRgw7I6n5
P4/ZZ5YLdvqprKWzbxSVf3Pk8Y+S5Q+7vq3hHl1PuHLuYk+Z1X8DC7Tst0/H3tvw
HFey0klpFkrIroSmyMMrDbuHIZTbP7XW2X3oYXJpVhC5y1UsbwoRXqn/caae/bNu
JDQiDyIikSW/h5KGPI5D38NWG1PsaYQcyDl1gVYosfQdOxt3PzW4aOfxnJ/x4RDQ
7tR77DzX2nnt8DgLDiDECepUvnzZ7SatmQb+VxbZ89ou9i0TeBxtHZZNkQpfkqRE
R6pMPACMQFOMso57RflC5oM/eJac+MXzQp6Ta6nASaxhdLxZkD6h7FAr9+4nFNqP
oameCpe2+vHuEUy2iplJdU+IgayoB5ADY0Nmo1JEc+B/ALXkgn+zk+TDeIo7nvhB
eS1olrAXDy6UGDoRfQg+xf0KFsK4j0SOod7ZnuHiEKrAG/UdyGhS/UlEgX1NWLzY
5/xhB+luuu93ffwlQU3K9O9s5f/ZdkLglKJAr81Yodj3uN7JtDHMctGIroOyvCHG
onpxtZHhXCtQT1bqCSFFug9/tP664upUZC8DyeDjrlN6ApT+yIXwOa/YW3+p+phq
bxmtN6koPFXeSm9yOPPyAoncl5u/mc1xMb2J6NzhyPdvkePTPsP3bLs4TUWQ1FTi
3kj62a/zJSP7r+fqYGcfODIRvx4zQIpC2EtWlXp0/5Bi9edHIr4repnda8NK/FeN
nZxB/cOGw1gACnae2lJRuRf9SABe28xuOGuFionvv+G0FI1QU0w1KiEXwnrjdHcv
XMZU02GPvJuiANVIiVvBlYBt2xMQXVgVwzOCCWdVi2T5n62F56gJ8Ntut/0PwW91
WK+dbm+jNbAhNf6eLhkQXnMWAHjCBIM1obQyp/qUcPnP4ZUDJT8NuAPVrjHEcnkU
htoUEwsk+9b4QVXuYyLkcMYpUnsfvYgszpl00J0NhmiOeh8yC3O8RSfKOZ9ZiZaG
n+2HmxlrB+0rP9MWZViYP3g/OOHqnC6Sy2SKPTnEPll62041qtUxXinj/jJzuKLQ
bd/6LMkHCV2V74s/6ochD9xu5IBpE/zM+8qEBG+jcDIiNgc8vDyWz4ZahXYFtZSi
RLFOLf/H7duPDJZDfCAP7wnlXCIx1s6A8/tanTPp/oMiYnM2aZnW/g5DgytmtUVV
F1ECym4KiMHtr3Hj8Ek5WfbOdWKXBjIDmhkJOM5M7RQ8ywZiVk9y63E3jH2lNRqe
pN4OnLy9UrkmpopN1JZ3v6ON4EXiHEIn1Qls/lkvTR+Ln0SDq4SLQBwsdvKMpERa
iKDnk+uC9re0ORlsrL1Vdekuy/10/NRv/Sie7vCqKyMbjTv1heVkIOnL7jKpWHF6
gVsO+N34n7oAGsMZrXJ28/bZuVEGpGfkuZzhN34TN3K734/SrPs8gf5JVmxHF5q2
KaNSQLXhrEsuaEI/mWhuODj34mkRK0grA9mTJex11FFWIaOTCEWqSZlGTsHX5vm8
ryl8oqSjnPUjruiV9UvbF7cO0a11+LYcwQL+KXjp3F3FJ+1J2mIyTiRR5iG8hjoP
PXiXaSYYwrxr70z4SmHd5jVX0ktndqwgUn2U4KLfi+IKCJysRSu1td4HgQbRQ/PO
HkoVUPd6Ea0bza1BwS1rXkekgbJg7mKxfCz/BN2l7PN1Wge6mwJ4A4tiWR9lSzCJ
gTkOZK5Py62hrtZvew3pG3AE5t5UXqFqtXC5qWv4mu3tp6VhiGQMpTBhvpocDx6J
odk0KraZzxoWY+kps+AuPMkqvVXiUdZLjWh8q/2KQQiuTUMr1x+CLkvd4sg8v9aO
fSW2xdEK2Nfa+Dn0yxYvFz0oijBbwKJjBM+3JiDey9xfbpLb90iRIk+nnXjJ+TwD
zF/1A3GPBSrlVQsmyH0/lAeI5tLCRXpnYz55YJGamZwiP6a9VVPm3DnhL7QsPz/r
lgluJFwWDiO2mmAfqeW4/2K/cA13F/b00dYRV+IRPhCgkfGFvxQhGSHTCqUVmJj1
/6pVwWeg8JWFZ0cBMJH6NWQQW84kDckWySdMjqOLPwYoQ99L5Zj2w4DUU3Vkx99B
KhppRARz51OEvP85fShbK86+WoRxBNcCAQUyhyuabeDrNUX1dMwkDsT20GCHkSst
nOl1UjxJPJdMNud4eheEKUIIPL6ENZolJNmYovAoJchhwoPNkTd7PLMlWXKcEggA
VMrqDg3EfGAjoK3Cs7wBE9WMQJP+3CVbFvZtxA11sldPEBWYzvyuxXvNvP77NnrN
z87wrntwlJmsfp+FMPEltRmksI0+m/S6KyLp6PB34ReOd0Hp4rlAdneQYerNdGyj
6VGvJFNmAF5RKkh7Qip4Y7H4Hycy4VnkXGkyS5A0PWv3WNNmSWgXhqw70r/UiDvG
nW4bwfRy6udjoTOSiE/XSOhWO0/cbHMqmBiRyJnWtppiu7nBG6/WRJb4iExbWC2h
Fq+tSw8lT/wMHvlz7lMkmhBd26ArU6NvJ9q/cwOk1vE819G7Kr/MtC6e2TxrIagm
Nc4exKm6xiM3+2lPNDlpghmtAAHg/fUxnjJwsoCq+9sF+ItTme45SXGkch+VKZ/Y
VRKoxN/dIpk3OUs36s1oR2fU01NDrUSUZ0Ckdq6GSvWL768Lkw70bjGH1i2CQdVF
`pragma protect end_protected
