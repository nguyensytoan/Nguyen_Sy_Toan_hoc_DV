// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
E7p6Ot3/aNVxLlAJOvAPA8GTDN6onKDRFeiXA/zjJj+ySz+ZlCWaRUFr7WtbvRBP99DYJfbsKI/1
0ZP0PnijMKjt6Vxi7x89S6ZASQBLSJy1UyYyhwXc41W5aTxhMGsAEaz3uAXtAbAXAf+4dRx/k2d3
ZiQFdMF/3QV40kfJDZdPwU1uh+6/Nr7t8BayAHgHaWAPLP3VkHb1g/Qs99EuGnCBNjtO1mnZFk2G
Gw8OT/UXNbPFCwYkuHBZYXoWFRk+SCsYdy4jV8kz48eTOzquJaV5ea4Ki8VaUpqmG7Es0De0zeGZ
Qo1EozRkBRdUab1TFP57aXBQT/Kqqg86eUvFug==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10896)
J9+sDpV0JB1d6B53ACPLb+xAHgVQeeKFqmEyfVe9GCDxqYUnc6np7oTwxBIyKi8MbN9BzkhsfyBG
rQSBzyavZfZ8MPTR0zGXMCt+elPSu5Bqwl2XlIUikBtfoK0xr2LgEr3pnKJeiKnJNY/NDRnNUmuT
wsFfP1L9G52PIqBslqxP9SyO4q2Wr1BK3Sgg5YVf7avQ1tTi9Sxg4gHOqMqupXdmPl9gyaZ3KmBg
6vMVYAqFoJbR4qJEnQXKXgBmRCezV9gNyagBZqeG33iMhGwQKtvM96shm2xSxCJRp5Yw9pGk3rK2
UHuvyZ/C63aKaHnjHxYbq0qwOyJVFDLn/DFv9aT3DImiv1f0I18VCSk3jodE46mkhMtipfusslrP
EeyzuOwemnd1KrEPHLaj4ej7JASv+T3VgXQeqQIjNAKJu/aaQJh+d7PPX6GB2TszEDOQ6LpLb9M2
ucxG1mPAEamwHcJBk6Nx9c3XDkZFUyVVh/7VmYCntQJDDEMMmvknMS0uMUM1u2Svlt0EEJwm6syx
aHWzDpnKNh1ZHiq4MREXF7gOsSDeybWkpKCi0Et22PJvw5fcl60yvhyh4teyv+/EuJx82XMlgX86
mDb4SQQmCKu1zS5qLzopLkLf3+PpLeYsb7aNZh/GWQnrpiDkEswH78SZaMF7Iy1T4+mr20W6DNai
GT7hSaZ5XGW9zWpD0BdLtvVhgqseB9Lz8T8UP1vglkQ2onKvykEgM8FXDqvQni+rR9j+su+MAVnl
yacq8OqJWfrV+MB8vRZxV5kJ39oj/qkOIfC34QhJvvCa/D1TSFO1fcErdDhFmMUsW3rCiaOjSl/g
G8f4Y86sWmZfufLPWy/OP07IKF259DEb0F6rz00DDLywHQ0FxV/JkxLYTNNFbefb7WXO8yL4nPZo
ni1w1dgi/fz53Q39JuMqdwhDSLa++oRQbvufT39d6Z3qD3/6C/nqIJUr5SAvk/59WRe3tQ6lteMI
mMhfI4Si+eelQNArHFrSg7520xvyYSgOl1rklvjHDDke7B899mY18+Wc1VbPVjFTJnSd8eryz9WT
6jtxIQOVh+OIN/MRlc2b8XVV84k2NWjDCqnqJNqwx+ObxQ2fl0SWXPDpB9M4W8AqZDONgkbanNcU
7EUKxkCVQ3RY9jVdjdmIgZRw5x1mU/F6ei/s+gJXz3MMHM2UvEOGJReytvScUtX92oxAW7s/nfDl
wW6i8Yr+PkmKD7xLsFdYhnCL/cAGB9GqCDmi5R6xGLRXH2EEN0xOagOxZeNWgRSGOQxkP1DN0bUR
H7o2qtBGQP7xdFWTBKL+GHaGDmXNKFIuCC3k1u0EQS5oLaqEjSGry3bbiKqSJF1eZov8GItAQyCb
0JYTSyMgKBE9KgW+dvuF+kN8BUcxpcdd9J65u3jXsz1hOPmsLDDd6fEO4WjJy0QA6rf+yjzI+s9g
d8VvmoUF3DDOypPGCK3LiOUDCQZusZEVoZVonqGYE1znpq6BAEvXZIkDoexMh4aCeWejX9Jla7Pp
+bn0nhhCzmICXiO9seVzSzQeGkk2szqqnMNAcGQTnHmE77WwfunV7Gb/LQTMiCSQwhvKRlYsfz1I
42lp7lffA+s+t3sQpKxSV0egyDMwgfkSAsVKudD52gBOGMBM2mQlCCQ5emzS3gsbe3SUkt/GvKJ0
CB+oghbQCqqutMWytc0Le8MdoZHCzOhWbjNpV/1wnmZ2TiTdyO/g5tVGEQIwn6opfrHjBgbSPWDG
oW5mwVlJ1X3dgLM4mDPhN31/xoo/NPTEBOM9kyDgtouZhu5P/reVfNVrh9A6116Wau9aQlB362FF
h8BZQiga3MG/4taWTAMNXJ+yAkq8dPGg66v9Adv9BNwLK+zBRm7gnAKiDmDqji5GbIjX55gfH2fp
RcxfmqCWcjklztVw500DhSGr0A643GsPwbYRVEbTjFP7qGrlWnrcewoZEPOFoj+JEp6mbvlogDVH
TcbAN155YAGpnt+rYRIyoTQwmOZK86rhWIKmmITjJkzuH+OvrvE1oyrbkJ8URjXltbJ7uzO7i4ov
TCq6pHPboc5gfWrhDe/sCYGbUGpSjY2jq46orwlZwcBkxlUypNBIkTlQJg7H1LzKwi86Z7pTEklw
n1TaHsgiTTloz+ArqdJEkiOSIR8w9GoqBqy4MfRxq3FL8N0sJY+aHD9eHZWjPEOK/yTx6mnpYPrG
1HQu6FYAJSd08dUZRwKqVjWtcMxtY6dJSqcjUMmk83RAN1hLLIGpAz7fAUjZNnY79SqIbGR2YlAK
mVqqRoOIBIJMIzu3ztlQYOu/l2+9ffMOaqwjt/xabGdGTXHNjooI4OhU32eUOj5syQa8Yki6/Ul4
su97IoZTYsx/EdILMMfnY235nkCauhz9Wg437VhwW+z+2rLWKjZB2SimI4V6Ez45qWHQLdQARAZa
AvAZ2mk1yaFEX36aYs6IxxboH8ZdEP1qVuPRFJF0xXRJHfVpyTVrPHS+1PgTIuym2cMmTepsl8za
iEqOP/f1bN9+SxXjTo+sc6N+Ozy1bQBcaHeaETvRSglMYFabDwQ8Qwgir9NzxBnCmw42GtrHYUVE
aiHDDqFnZSsxiiNjqCM2fKJ/obmRLMpjj2WCR2tY+lX/328Duf5MLH2ED+6hE8eb2tL9Sars+ENJ
bn2MIbOlwK7pZGay6Kw/0DlTM00/t5YtoF43JAjhWiQaoaBfxGvp7LCwEqgEeof22eZvHSL30Xe8
FbEgiV6bRRJgyYMlIgcDt7VxVBVe25EWo9bdRj1vWU8osX1zn70qNA8P5Gd+tDLk4a+Wn/TSYfPW
v7yIu70vtGyaBlmVFq0MQNa8Zu+Sssx6Ym4MYcO/ExhRgj1NQZ0kMlD+aWscZ0DJ60fSe4YYrBX5
1oCcYDjpk9l3fVYmskbmbSJCSiPtd0sKy27pUqF33+h5F9b5/CdlvmLNc3/uiH3OqDsatZXCqD1D
cJRx/Qu2mUhBgWp0GyfnXvjoi9cb0FIhjfW80CtNsrtnbjBlF5tHgrudmDvFHXoLizptcNxgOIHE
lV0k62IBwF5WiSmZWQtXnJXcBgjOCYT7uPWTfajCsezzaowmrnLSn9+t52khcFSC4+lVefsd8Yi2
zUyNIgZ6YNb/9x7zovQvwkI2iidZF+4tOpVRjKSKoUahMprHJ86uVJh7bk6uQVWxGT64qLsoTGsv
hzmLK/13HfMkyvBxEAUohy5l+lv1yefqUvG/eA8Lkei+eOjs0jJcZPAQPlrj3DPLxHWTP8/1pF1d
kKhvxF/E7FZCRHPKbug+v8ggWU74YUEUk2WcDwCNgaQS95Ei0iJWZrPTTYEY4F3T4TfKOtc62VVK
S9hJQX6XatYsvs8ENJ86LzvEPrAx19tkYDYb02wGC5Y262cPdpEq7W1HxXLgUTm41UK9XJGRRyBA
wggXNvUokDjd4lJsT1p1+jngL/rGBkVxYr2rI2IMfkJFuiqlwbTmXKXbvB55EWNI5718k576I+gT
ZEJddiSVr+ZrLPbXkmNZFIDHy8uPtaWXEjh6iSwwyQB6z0Lp98RSmlXe+uCyKA3NSrDjLfQ61Ir3
4NfjPXBYNKV1hEJ3WXMLxJ9WjHI8IscGa82Z6qRLKzkSvmyFPyrTg1pmjELJNX47XWPv5C6DsMLA
fuG917UZOemgITtEL8uQrQb01fbRnhy8TsPNruyWawgngCBwwUQtFHNZneSamE0xGF4t+ty8idbn
ERJXgQFbUw9HKkJ74VrjO5vzQuvQV4LKEvNhCXQt/1q2eki3FZrXO9mhmP406e9wVp9KvYIGr2Du
2h+ptmHIPNKSSeZB9Is6SyP+2nhaa8QYk9tKqPJjHLqkMz29Cbg2aLbymwTbsysyAjTw3oHVBghA
ynU/Xj+wwDrWjRv9l6IjUhw5zWWcpnsnrNvUh7Rh1OxZP/jlphT6CZz34hSuy9S0LnGGBSeD7U12
fOonYUDhZuzwvrXUEHbosxZQwlefiqW9XJhywGQ4olGZinwSuYjMWxzyKR4nemzePrBtqLgVjy8Y
XmISmtjRO74dIzGxGTedCPThsPXr//dNBMLUIUxqr6sdh71H1cvpln1z6nBtfpIXgTy5PkNYOGaN
rgS3IB/WPmtFoir6WvREEZK4mJ0PhbYcUyffYW7St98KIgLK1ettzIurqL2g08tLh0DScEOHigm4
WbFfhhawwr1ScX1AU3/0jGLYIlZ6EOAkGycFQfFDFQ6sqCCUW/hzqxm76jjNAgC/LcLVqrruTzap
0Qfohyjv0iUmQnjn++lrjl3jDnyj8vkRq3ZynM4dz+gv/CeDKu5z9R5PCnnu6TEvYN+4cUbYaX+B
CMbVH753LuueyUzofAG0dneJd63txNWTzZiFReFXJjkpEVQlApvGOOwSNg8WTsuJmGcq2BbPXrAj
Tz57AX1TrSzrpB8vGB+WzckshGSCscyXHbsOWcoaDR/vHMMcMRvdvKgPHvjyNAq+cu/PW1QIUpj2
WTCgQ0a30R0E1xGabtNvHbPBEKeYoxnXoKLFLgBQcnRJDZsieEwMu8Jy85Kj3515U4I9pWYIiclI
p+Uoz1lkgXyQvsqNnv7bZIkBnCFvhcBHIfdiYEGQsK+nEJMOdSzge2SLqxnwK+qGire+DB0+386E
zk9Lih/Yv01OC13EUzr3Ejahrmn7XHuLsm2j4QgWLJQJhPPDBlMflezTeRr6MFyOu5tUUDhFB/xd
BEhbsIwzJesftD8pDtZKBYO9aT8rdL4nqHDm2u7/aEqcMre1gcXnhpjZQ/Z6NNuiP3j4/PjmyreC
dHqYW1pDneme9kYOfXfsG7F4sIzpmmx2r8SjaYSuByljiNM3HcmQre2T1eY0cPJDGCDVN1a4BjYK
Bhb5U+IvuB7s+F7zULTvYCgrA01MMxRAonqaua/bQjUhI2XLZb+XgViz3/uYdNFthmxVL1x2urA9
0k4/iRjZd93ItD/dTTIuXXp4PR5qJ4RhqqvyaeYY5leUSO2Sotdcdm/h4lSAe7u5OrwDAAbhJ+Bv
zZlmk8wcbZaT9dzvGr5E/m73UnOxcBTHueok/tbn8Tc0hukh8mdRvSv2MhAaxaQmwMT1VPByGNHe
kbX7XbKETv95+zKLSD9XJVnpgVdoL7iNs69r+d6ul69CfvzObz8k63pppfxnmoAcHYP7QZVEj/Md
lv8ZnvhAk6nqJULNHtdiZIISLLCxj+islv1Fjbjf7l2IzjVA6iPdmpKfdqs8ZZfZWEcSsxcdVvZ8
n4J8eO0tiZVPWJzQcbaBxgtSwUK9e6meNcLNrgZmhMo13EaAW4ZNCdOLpmPhyevRpleVAQQOGZhK
MIAf3RqQ68fLV5bcpQPrdGOs+Qzn5vf3uBTHscvhEGKI5z893hF5Uc1XhAxUVlqlr25+otyQOVUn
08nNGpexx7p06Jb7602l/ePePLAGU4o8P7fcuFZzmbjzsDoQcOu6Bl9YfZ+iAvH+GsrLN4CBkz9o
XYw7mXdzkxZGkbEGxG+QcmsCYcZF768CkyKe3Qi9rtl+OutzhMq40ZoPSmeUeACNZ9LN393U4Jtf
YN1F28N+3cYb5PXbCAxrFGZOH6OxxeF21emiFK/mbn6fanh5Uw9gZkBxco3pVmdnBt36dcOswi3A
2jKiM/JvYQIR+bXWGF5a6fsev8AIixdJj/503QR4zHPECmlYMeTAqPc9NT42ACQ6I7dT18JfXhZI
40RE5lNvGaYGQ9gSR/Bwt4i7LUiQ2m9DZvXnBM3gOnBhUDmmkGrYGh7+q1fTuBwZpBo9cU9Y4bw4
2AuA704w0t/vIwIAaUWwhk0QW2xtKnn0hZCIgNO94V6DmGzWwJPuyfZ4dIsObxY9rsougZUUodFJ
p415CL7qFrZbG29sHNYkrmc+nszMC79TUZ5IVzI6ABhww9iBIc84qPKyHEoOKQDlPN9OVCHWNCii
BeLX8VH87kqySpPQlyOVkSwbjjBqfiJWYrgYLO4UvUqATItWEN19RPPJt0Bk5sAhEe/XhFpz+ptv
qx0lMqV7tOy5XaE4IK4MJ7vCzOQLhGiRjAnOWUw7KjsNWhr4P9l2N54zkjMCHT1dv7ie5/fpGk0x
e6+skS3eLiACWkioHVDDEmRF53HWxfwa5977ilx6OXoRcNlKLT/vGabzZ7O0fSk1n3Q//r7f5e5d
tzKT61Ll348MWTvM2GGBl4MEp6wjqwOk+g0wyt/P7nFMhI/p80pKci+J0Hj8g9LiIZWYI9PXWa0D
HmsY892ZEVb3pNt2zXdvAU29lPvDIs5pBFX9o3xY/EwcfE6aO2b+Hzh3f5dhhRoDDL3lWebY9aIV
o1a1aklA4NrasxCs/ondsc7J98bPQIdKGvveIL05Q92HPN8CJZrAAK4FOcLUFPnw1o43KnlNjRAF
RvrRrLvigM5/yxLhBY9nA4YBzAcs2TcxpMLYhkhN/sjNPeWOLb6PABVI1tuhTDl/9xiWYVlvjng1
G4GiHoJT0xKRdKNK8i0JsPEfeK9upmLJAGNrROr7IdayGvecLNR35UZK2KtKfigoZp3r08ezu+Bc
KgBLhwDDCXu7zskKyPXpxsdq2jmyDHGa5Bh/j7fiaiaQFwqc9NKgyallya4h6UShWhrsX4EsTK36
XFdro9ysE0HrkePiLo21RGXqlktbzbGAjfoqXhPr2lSH1efbONcA01C4vJE7d6O/T8xTzq3tSH4h
F8kxb46IvO8lDuR/HD9HdHwY+yS6RapPTUW5WwuCZcLIixeoh1a4hd4bOgRrpRY0jMl3f4vK/nwo
Uuz4Tjl2w46yCanoKWFzlKR7B8bPg3QYUuQT5Wgnj4aVC5eZ5S0+CdhDuTv+dsLD11yCKUGage5L
cus01qFKUN+gegknii7VtDE+IJ+9+uzlQab/7skyHemHrG+SYhBE3MU/DXz3ST7S5ZgG9qjABrNa
Hx4utTrw3qXk28JPj3abaLeKlS4H0eh3bwHlrfiV8E3emU3LqViplexLqz4dmEjHDHxtdYY10vqt
akX44d9weYwnS4KSYpdaHohj8aaKqP2N+GdLag/aZJUW8OLXs4Do+t5LPUI6m1FP1tVYErsp3KLO
aEPnUyQqE+m3tbqnZghI4ZqsGLYwzzg92p0KrF0vPSPkbqGKcZigI/zEfISXG20CD2bGlH+Da91F
HsyhOEMeMVHHpprnOnWAlXmragxlVv8zjnzjrAZCgUFjKNTeFHp8qsliPs+DT/uf8dtki8P7ljnt
qn3bikc3mKIANh2h1YDxpnjiEkBybXaEOteyC2KLekKuknVFT8jzT2IKUv0pFrMIyubKjf94dkY/
Jo21YCpg/MxJ565LY92KkYZwEE+uE7aEb9b+k90JizNWD6ujn0iJWL0DmL40afrNJgKSW1bb14zD
j69FNRqaKjuWwzXVC+iUxhqv0z23W75Ic2Bk3D6gzmDJg04pnL8uPCDLFTe95+vZAnWRNmsrYPcF
hJvRS56+Joy1di8MDAeWOz11JCPqVIPoAJiCBcMDfPcxW/ltfLlDBlu8h6T4qlSKJq0F4NCJX9Wg
mV2tV15HROiC7HqzndiZXEBSlQGWwUDllBv3+rC2RIRCzpUMOL7W7vVltU8tlPQIfeR3pbLFComU
QBvw8s2kwMoLf53GOmIwXqD8FKIynu+z7JRzLn6561Ai+MVexexOkmKzYeFnMDBEl7/LkobJLAo8
xTy2yVIIIwakEub0hAHgacnEr6IkkHgtLXhg5P95iOb7wVjXZk43/ahz4lkuX/1Uu9N5l7ejNI7i
JdxJh+EL/aY/o3Pe6aIrmQvenuiwBbpL2GR0c+FypHcfa1/gIAw+Mekto/xgZFU3XA0sUs1aUYqe
pPIlELOjyTVFYKTLmxW6LE57s9aT9DWKdAQvO6ZaU/JzMMJC9t69Di5x/FK4t5ebWIEm5AjnQRCq
fPgHmxkugRPjs66VcsbOlMv48L9ZAuBMLRCGlo2VJLGE1W6kvSaX1O18Hk4m8Cpuw3p1huuOEUGT
7iidXRezIz/1uk1VgBZOF1rjb4y7Lm/RzAHNXKjyLYlYh7bK+sQj2HJArBTFcndA0faGbl32vEZf
utCpDI9Iv3sGgRGFgnamv62YXMQuk4eNpqrEkG7ojU4WqWOSAhylAIA+fnIGJRi9hc/UEyNbiNy+
DFxONMi6Tc6XHwQEd0UVyhrdSBMPbmvVgHVwf1zsOeBfVWimQyZBUHGUgAZc9/P5/91xqndFZC+u
q0HTlmCXdBqAgMN6LohoiLZWOH8IbeWTOMG9iHngk9Ivcv+IZLOu+eBDaKh4xmCq2+PE2NLhrG9f
a/WlrAYxu8Cu89hdVzZ1bTvJybT+mC9JM1EFCLhLGZPFrFepBrdDqJqLuItcG1OFLclTWr4WuNpP
Sz0oxSu0jtayLQiq0fFZZ+/qgUdKaHWEeans6gMBE+QXaRLgkL/SSGfWKb0gSEScGAPfbYeQtruq
T1GWqSS3FKNBZAMHnh4EJs3iTcnPf1ohsmiYcCfD4JECRi7On6JGGrS1FEZr+qzEPpolNs7QumVe
VvGM5uR+bDXd4OmYXVFgHHxVEi9xMG89BWV+gzqMcAb44s2xHQPmg58Vbf4FEeMkiwGGmvPBc8J1
eNZc7lo3W7J38pqRFWXrQD/Qr2SUy4XEn67Jbm9/qMtYtya++3QkTIK9+rPNCrcPjJt/LWWb+nkj
22Kk54A9gQCpbo7AM01buONcbqw6QYFoICOUaZcQKgHIQ81X9/LlsLExqNc7R7blsokHyn1j/mgv
oT22j6GqOVqh4TOSHC4c+0iql4hLDPp/ZsXKLllspsf/4d0QWTjw4BXfaaVzaHZmC8GWey6hSNuV
wZlEfTKQB4gOdUB1Gfk9H6ot9qLLAkX6hMjB90vUvsYcQfB26VMR6AWYsQgYL+0CY+tAESqnjPu1
fUdH4LcOalX6hEAlYblPg2ThNSXD7WDoQzw3htdJxuWMpCS1hJE6FwrJddVujb2kPaT5HV+Fm0bb
R4Dd+0KR9s6KUyaqa8LUMQi+gpqkNpMfw6P8686GQZzhCnNz/uB1JIJ0Jf36y5dWZUxLnrUwLnlp
Iq4eqL3/dP8tiWbySsmID95qWAWw2vnIeqLx7HDOfJL3kEAsvjrNXr/vORsXeWKJDv3m995cF77p
2Ln13XtCC2ecSjbLQIdpqdiEJHjQYgl7cnGH6fm0w8wmdb6X+KlIgMr/v6l3ocOqHzHZskEy+x4l
z/CAM5McQ/XaoFcor9oLeCux5g0FR8SBSsTa9NrGfjVWRK+/tbGOXcX94Zr9gpWcy9Orsq/0CfS9
ldli5oZSTIKYgmH68aSl+OFsg00txAiTSobK5RXDwEp9gs0yYzPq1DqijwIx9L2ZUk9bojpDH+z/
KwZOiEWegtXru4wAKLWgYXJogYrZnLDX+5m22DAPm11HxHzreHpX0qbKLRxnOhIhPb/d3SZLQa62
SFZEV75TlMiZv1Q41orPRBPViqyzIuq0f0hA0EoDwFRt0D7bZHbq4arpbJxZMZymosD8HAV6k+VF
BFzqpKEHuetRbjYcBcOitRewG+0b1nL7cIBx1aswEKdgvdPSDD2Ps3YZSFdGtzRtTlkCsOI8Hefs
V/7TwHAXxYSjkXMPJ5PgoDTr81sNS1ScS9QHUpN9K77ZQ7VhC6XGOvdt4AVppfUxBScGfdtmBIYR
eNIqhIpfdYVbKY9LcVh6TEXfWb619UVgbBd41z0TJLwQ0rpzd+Y89adEFTOiFeXRwGoW/qO5epGx
d97po1tcpVvCar6G3JmFA5TnRAWyz3I6zlIgqoIeP2dKF+uyDjUCsCJiqZdDTwEb4fPpEU3uWW+L
z9kTbLrAhjeDrQUqlIkw45inrAku3Ltg9FH9DEXKM8UUYfQcB/PR3DoPKefe76xz/IqmZH4b9YA6
GsBj3V0OuRv18/i4/cr35UZjKNd9GWPUS213piuLMhqiyZCqheufIq8F5ptFfPZCEKNC3UO7AMDG
UqLRwFWrr/XPEjCXTmDE0Uw1ylCqdntNZKNH0fW1LvkljdKZBNrVcMGjpnRMl5ysdYQiDWlxouFx
K42RyE1pe+AMMm92tIhU1A321qS37UOz1/ll8dlXSysTLEGe2Cq96AAlfOwGHj5awT9K61myA/tc
RnirLm81d3m2kr2pv9feZE7SzeD9qg2XE2svuNT8gQu7XRBM4rFw6Fph5iU2zTr+/HN7SVbEJYJi
1GbnPO+99D7aZiWo2i9QHsldBgcSsnSCMn2BrIN4SL8UryKeh/gpPlakvXcXlb12ZQ6hC7EjwPZW
Tf1cEzeiSRPgTGaX+HOjSRYtONJ7hBWnfWlCLcLFv0QH0T3t53esH7/LxtzLEzxTdPL+LP0FMBDE
g/tQgOfWnO6DJdV7jpmvB4mVjTvHDaC/JfjIjRz5GJ8Y9cREtEK+qF2wU6KnRUu0mgPJbHHUiBqr
GyIcud4n5KUMRHVq88ffWaMtDW/WSzMdDDeAGrKj/B/i75c+856C3EkGdIOZJQDjjNsont8i6Izc
v2HiwNE2Mzz4HeTyRtcL3/ddJqTIZ0mL0DeeDMIdb/QJj5eQXJ3LbWyfMsPeAXkBF3pLGEE/xNGq
aSS3wlmgl8hrv/+vWi5foeka21t3VkacxZqAFGcW5HiPgiHnEA/htaS9cFqproNR8GtQBmLYJ7jK
EzVUl2zP388m0t21XwzYGfg/U4TH7uuJPhNaNK+b5cj3bnpaxpYdVhS1SR6GmTTsikDfJUxlpdfD
znb3kN+6PGaaeiLxEGxnds1CX1e5TnjdWc2TcrfYNO4dp+gJORbyVZN4rRncgTj5Mx91n8bRfzhG
s6DR1AI4DKugtVAJ0ZpA4lgLeIWyxiN67N0Qwa3u7H2n0h25XBLyE8kxli5X9zeN1MP7tXJ+94+U
xBb18beSrNlRVroOOC+RMa7MDuzXq1KCPS2pGwtqoU6qNgBEtJgWv1mhqvCaR3K33gYgYA33kbEx
4GPAjvCNzHk801jXcZkubgB03es6mlqFQJ63zJ+eoNiCZYm5EsNjjMt7TBgxh+pWYEwyZ2xTWKHH
Kx6izQxUue3AuY9hp103DADNFqrszhcdtgaOIpaOee6FhvVqP9DDVSXov8ow2IHyqxk/z9lEtylR
yUecoP5Biw/PQOJDqob4l3ZJf1rHo87wA+WWqpuvMdKxG2l+5cuQN01Y9JgMfngKD4uFi0WhcH2k
PzSSrhxdRobB+6M89CGxSCyDddtb492+xpJDzzfZrdokzLmR70PT6RmJigR7VETTTLUd23zVZi/+
xtpRWOkK642Z5G8suJGpQkGw3pUHcusRtGBP7R1lqO6V1aKtRMUPctw09Jf8K0SYXedvFKPREOCI
uI4thzCrhPX1qxNOt/GkJsUehU62xYmxhktOkwQEBuVZi3aUlJDAMOYqrKAz8/bCMrg4GqifSVyF
ejt+7WfSwAWN44JrdxY5Yo0kzuh0Mdb9v+3XMPJdzmBUjaafqzTsC81d59On5RjBfBOCPGk1xy66
szGdR+akscijSJvvnDjVfLzyf46hYlGBBtCNzvQ4E0DXLEEHjHycZDnDXO9DzQEjWELbEW+tLzWL
cW8fgZLZUNOROExf7WUBNRV2nNvbN7ba6X5cDiwMA/tBolZRTZ+0xJx6JCbK4+Pr6DmQg4ztD0Tr
iBYiM4UoJZ8lZwK1aXJsE+X18eRZPLhZFzbcN2KBpLMq8HIuHRVlnX6YZHWmpcVTavvgi/f/jkyx
BzSwu40vv7HrXh0TRW1YRwWicdLbBKviovuNXYeR/VLXlzOZOojA9NLUl3BGzqcaZtmPzQNZPO7S
iUlS8YnbTApXNe6crkPaqgbqi6m15lkyUCgr2JbKpd4lQAg4kkyPImERAsWxT2sHUFEz//HgPNOv
08vGU66RJIAdOGtOMWGZyHI8xFFWHOxjekwMT+EwJtCUHMcKJOn69gdnTcUgxbiCElM1hE5YKBC5
BfmGGGuWq7+5sBEcW8i/urVDie8/7x0Xw+dd0MYbKaNr2Tw79S4i/5FS1U0XCIiLwvUsDtifyX30
5U/u8H7O5XZftMcSJ9hGYO+TkrIp3WSZHv8t7lV6jTqZiXmg+BMOz8UFNfEbpJG9G/1TOZGyDgVB
YPEt4+07md4dQ1Ih8ga/VEU7xE3tw7KXij22CIdc69jh/60W8K3D6/RWQ0WEKiPhyf6v4mi72WZC
8/xjbJ/YwlLEIORV5X+uDeYk5Ssu+gLbKxj0Bab5jqVEEf2opOsoeRCl0BOFoA0siOdKl4yyKx65
T6aTSFXHv/qbL8Sz9iPk4SYchYsKrFtvxeG77RXytV8gwJlxaQcSaU7jepbKUxtqEN+faw0Yg4gt
jOYrVKeVsn0/3tkQQ5J635d7rUJFaGfnQ8Fbw2qocR2KoLzTM8AFFHo376Mku/K/les5qG8FDKrb
pSPYqki04g5m5OCpdHJaIwpUmCgCSF3iSICtAzfMIty7w0HHGTpPYDHG7IKrrHgbmgb90BqUt67b
Pb5FejxY17rB7y3Y9G9ncIyTXGkfIpMaTfFMrbCpqC0avboDS+ACPxyW7Fz4eKQ8w0c/QPEHYtaY
9OTdmgN2Yejotvx+ROEkucDcu+3YDa9vEMBk3f3Ru+Cs4ckTeGSlPJQmUAY899z9ENUL1etnD22M
SaUFGuFFRVAkLqSPrlfn/oNWY3KEm5o4PCLJV/ab8XeeSZYbK+S1bRlIn0ZOM3h3WK5g7OgaAwp2
cVl8Xl5v4njKilNy9BydDCovIIpxidLK3MsYfLB2vCJgoV+SGUjz2vyrmwCIMd0YCxrLZ7QWQuhY
eA+nhrbfl3t6qOGVS008ZLKgcK1yjbi067u5GtRNMRpbzR/lW7FxbAI1+JXNOijQPuU85lzVwrfj
1bAOEgMaQ0M+vnMSqy4zyXlqApbvyug7jlbGjPJJKTCcLalEGsbr8gaz1zPnSPTco+t8FNpWW3IU
oerHUpchdYMfU3imWO4nrTqffKUfm6ZC4/dFV2z9GkGIxeo1H9ADzXARr02BtelNarZwUEs3mQ5/
UAiD2dMoaIfy2qyKiZjcwejvhCTRfcawU+zNctnWhWKjw8y7LFkuZpqiRI/2rXUpBNlLreCbdFSl
gPZ7ZZ8Ur/kCrWO1m8QP7PsVHMAQ/DZ8Z44j3f5p2XdKn3PrmDfyx0b2xtkJT5q40NcvEIzojSbF
tHFlNIv5wQ6zmi1YQ1MQRWNNOCGjdxL7TfIrc6v+cuFotvCIL5GWQPxsoRuGDcLRfCdcib6XG/oa
DWm3Ma3kQa9OHSC5bhr5fMxPj/plCGUn893x0w/bnFO+9vX96vF5HXAC41eyAhPLEvKPJvCcT3Uf
Jh3Uu+cDJQbnAkgeLFaluagHqdWIeQVSwEAmsKBtQZ5fYNwhVcm1g/E8+zELjEEyI17vwV5hf5mU
IuD86xByaNpy8BsjHfn2QEOSl/vnVECFkpWpvm08dXs//yXj83sABPhnF4iacOtdlXtijxZLo2Dr
bfgTyfjIvBjSTuhlu6X8cVyes+Po2OpaFAQf5ZgqkwPi3rSfxoOZDsXgbFewBtw3PuxL5WDDcl36
i5sViZU+A9QhLeqHVnclJ9q0jTi/11EPm6obKanoFUuJhRxPzmhrZA2Q4NqnfNyPRIO2eixhJaMm
xQFZ1jS+JxKgWfW5OVhi8S8fNjpAC17ZiZbZUBAFLjrXWzw4ysqARqlvqmACelwDxkD3IkdB9SeC
jUDjMbJTGpfwXG7RBWmdrT+B8XhnFoo7yoLuxx2BLDo5LFoM8I+Cpl+0hiJUQuf7KEo9bqOps2Xw
A0YaB1aJ3FD2ogjOvnpzxR0BORsYfjF6wksNYJFErU17WNP1xc8M/ngRImXTeAAPRU4v5u/p3gXt
ZljYb2N5mTqIDHiF3FyfkFTC2ihZWe7Z1b+YEVEXy7lhUHuAwqfvkvF6V51A5wL6A51q+sEIIdOV
qDBp2fW+CPW7doQyQxB9hMJPri4NHH09iVKqVUQRmWXlzlewLJyEWLaehGu6qFu9ltehWO1PLa1+
aNAPt8+ZwKno5/y66kIy6clCGSwH+hL0Hhb5fr65ZDe1b3bE4Dd/MlutAXUs8WWqyy39ziIb/FNw
0lN4WmlptL4t8oAzMlMmNxxEB2M27QNy6zc79zbT0lDOdBOcu7020cTZ6TxbYfzh7DuLtrSp2q0o
et+HF02krZ8GaxuQfGeQUSClRMUALGYfC3SA+v4x/mV+BgesUQyrSYiBqxjOG+HU6XcJcUNe2t3n
hrm2eHH4C4td2kQkwlLtg+uL7QTeUYbQ41Fw9ciMQgyqsus5cWn27wt3WeATbsLv0YbvKFojwtzi
dIl90k1iVb9S9REJW/P+VM5JIXmIwcr8VDYSC8RzoFMOYG5Gsq+doZdVz1/OZFGKUEn5zMgP/FP/
atf2RE/gadRwcaOxOjULrzzFsj57R28aiAVRhzDnQKXj5e6nC/EHKP0RzHFzmzcS95OVaqGw6LSP
UwMdxTSiLLJIFKNlCWlx3EDXJEJoa0dnS7+4mvqU7Czh6G346IYdDQuUAZRj39xXOz3eWrDjPh/u
cVO4s7lmnZi8
`pragma protect end_protected
