// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
yfFP8dEJlKCtjtFID4KpNA1zOxwcfN4NEDEf+9htLBnjC4LhCLw2tXPgYw/x9zqf4W/0ePNIrrf2
/eoRTypOf1f6fKiJsRrAt7C6WNEK8pGKF4dCVatvxDRI3IrkXJh+l7HSOegssZEaeLZIUIq+xp/a
6ivF9DxHKSooHtj/CHC6Ra3CTd4he7rMfj9hfLcj5PzIRoRp+coKPvdw+I2xd+vhIjIPXH2RXZTY
cSx1+J2c/yl49A/WWMzO/Wp6eRQePx9dnUBzqb5jPlFGwoVd4YupFA5See7r9XDvr/H/bRlbL11V
mUWxU9fuMSv3eRUcKMqK3kQmEYrK/2HIssOp9w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7184)
ccuv9pNmAH1sj3GnPSFpSu3WbPEt15P3Jz/ZfuSPz8PKvqlrLUtO6RyAbd/0RS1Xkx6kfdkh8MJe
E389UDuHRVoboFTIEf9vxfxP/w30Ep1bjdRdGl9LVn6vs0t0GaoMq7Z166FjQ8GeQLPbkhzqBrzB
7uqjgvqyW33xis7M5mtb6RUJFfv3MbqlXkYoFEThy1iMPqtaFzqfe9mtw81nrUS+4QTpZtqYpZzr
bn1Y2t4/qDq2Ml+AJIx10xc5LnNNgIucJ1wxEThVnEzsGkisnrUTzHka+gEGILtdQEVyJIcb0NPR
/QTVwZGlYuvV7k/MmPcjYzUhzSp4WqM2TXbacpBYfms8LKOIY9oAP7t7ZM4UJlAY+EaGJByv2eij
KAw14qIKp63spLmrf4b9viL63VJSmBM2F9aE+m3lATuGFmjac+JAg7o9BTTbIeAANXm3frpFSNzy
IG5jGb7qCKKbm86pQWg+bg4yWBkMa8W4Zov9jhvxUJUqf/7HGl3yLcgk35wk+4/IsVVlXf5HMaGF
wUHHZA1alkSVQiPkKPMZ6o4bHY46Eq0V7MzsL5788AbRktluY/lMFRcoaOOz/OMQlsqGrPNMcplV
/Gc+LVfON9GVrmbJD6EebsdbDn5r7/B/lr8bkl7JAOOT3pDXvcKr0c38aMVfXiKacq+I8JdnCVQ2
dASxDQyo+jBx6yCHtlD14Wr5pjMXvhD2anj73aK9GG5pDViqClWytD9FkM+lYGkgeKyGA01Zm6lO
7LC7lgMUIp1kbLW5PB+5WUFi1jnmNA+/1v2So2e42pqCteewJv7IUmVLD5OsowNMtp8755ZMlyD+
nDdE9pxUGAIwTPDYbHriyK8i49fR8cMqz8LGasN0svFEJZcbsC+cVKVSWeORMGLAiU7BzajHUYxB
18JmW8ZvVzImCwEy1Vl7YIXZnciiS9t1ZWmkUqdwQ8XUoRsF7JHUEiUA5LoH3mmMxu/aXai6YvFA
5XfJS2NEUig5mYdYYKIxH3lPITSLgi2QwJyFbyIBIL7lR597d1MXPHpvVrV5OBUSg6BlWIsLzMbJ
uEtJ+lJt1vfJHf/ElQ5YYULcvEMOpkyhAtJ6mixzuu5ZmBiYVsSXrt8sXVI4H6mJqmmGiFelhHq0
yt4oXG8m/NcjRGupXzVCaQqqBh2YiLyKPABfkcR8N4cbPz0ajHAT7USx9eukFKiv5zwrIaJWQ1YE
tAe0eoaSd35o44QDfAEveUXvGHpWvz7lfB5p03HE006lUPoGz5UXRo+Uqd1/ibcnbjr9vccPzKUS
tHYskjuv0S14UYSMYwMr8JD7PtCwTof1koFciXDUqASanA5/ZdjONxS/uDrkdLS8LS3EIYP0TPEN
YNmP93BKd37Iy36u5d8l/wMT/Lg/UN9X8lIy36PnkFb5TJsjB2AbQwtvusx19qijCsFXqMlLuUEu
otBzd5zpL66V3p9UvwodNpsAkN51UEdoxgnNHxZ16MimT9tKEb++DbB9QljlgrvJNG1U2jz2ITiD
Z8kd2vQ0rxtbset8pZZSWDSTwJBPQtqacaTu8PH3VC62yvtsu3NZ6hv2tEazW4P0H2bhZNsDk8eA
dnJaapXxfcVUm0SHCtUpXMmT3Ah/bXwpBLI0iBwYQ+tUC24WCi4/8si0iji0CyG9T/P9Zf7cXFEB
KhuDrD9l/MW+v4+7ign6dxX/2+mqwatRP7RAu68prsADUnYzX/Jvx+QTFG4b6SILWejdcOTzH8Js
ZqmTqMQd2+tajH2KRWFGAdLp7BgK1DhT6Mxq3T0tLg8bRVE6tvqdVrUXDwHH43ygFB+ZqWWX7chN
rw9rFzG+pLer43vsjn9E2TBiWoqiywwLvWyENRzX0hY8SBNKlLHREZ6qnxvMPWHMB+xCSUht1RIM
wS5qFoH0dfrufmS2WzAg6untbpgJtbCr4yHguJ00tfe4LLt6IlKZfiacdqfuke77sBN6STqPTTHD
SbJuPGdyW81H9GnXpUG1AA5THTFr1Ah7mZ0PIpftZK7oPmyOyNs/xXcG6WKFvQXRU6Yf8hZZMlpq
ZHykr8k3HfAHSxUufVhhng7JaO/qHjxARrvhWTFtFkKDzIQpiiItDokMZHgdc32WtqXBI8DJm/9m
6X0LrUBk8V/H0Lq6LgKw5no9gUwchAO2Tc9i93b8+ZzYEc/cA9Ebme10/LaV/Y60phES9cvNGbEH
HGw4Vq1DYyFtrZlHyAYlX5PaQ6cyIL+gMu/cpqokbzYJQBCXnzt/RlGDgzi4wxPv4m/XGgpr//2V
Y96/YuOjzira/icwwdH5MTapFABOjykrRhCZuNuetBbX3BcGLIdk7d3GZjchGXKeXCyyKtSw9f6v
PqB1YuhybsnuaYJgAuRtdECmoJVQMsLb2AjTEZfHOCWoRPgrL4k4vnYU/7XLHUisJR3YUSuTLpd6
OJT10/0+nxGfNMjO5OLAKQZbKsFdnHSOkq4UD7NWJyweZig2FYTHhk3B44P+8P5v/ES2da2QVFuy
TMan0T0Tx0lK5hwaJgjN238PJRmTAS0W4OdPqXcZAjCe0jbojVgDExLewQind/jiFrDzg5bL0Xg8
5ZVed3CdqYsDuYWUb8a7Kpu05OFQSREPkgTcCSQjs//Lhd+eoLuWdzOeYNea3qGs14dy1J/sKYmf
DEwXQkdh4nnH8QNEsi8fbuL9OV4oLEhPuJprhCHQeyzzu/Z8lfX6uq4PKFfscvR28KK/Rgb3RIhn
Ims91Lv4B2BMBVqySPqDr5u1L79EqAO4adhxi9OKAiXj1i197R9GSKx/5iGBfbSiCM5uYMuaPCjB
2UqF3FKlma1l8T18dK5YNRRsmPqhR81i9PPVfvDv0xFIwqZRKcUat/Xt+eNJvexBkNWZOGVUeEi4
29DYs/lXYQrdVDqc2iCCiGl1pNY92rBNUzSGZ7PMaEbdBHDeaNt3zjiln/O5gGRLsqbAqwb+qP4G
6+58KukcdprdZHDmMS7CMaWuMZjJqRFC+ziZlkfIqscaMtU7Yq32Hxi1fJuRPt9P83HOJ15CEMig
R4kwMBPK6E9swdmu0UJgf54lXXKCEY+41RJ4WbyxibieorWqpEFkiVA4oQmcHq4EBPRPpMThbsu1
jRZhip4pVq1LbapOoN3L5Qu2pR2nHYv8F4YuiaHLO8vsiX7fJoyoeGOczRPX7i9p1d2eLTjpgc7T
hEEpSt+JtilrPOSV52hCtrKY7zXzNVfG7xc+OeHYfBUVFPbUAVNMn3sDNJ9fe1SO66ZhJ3GrL1V1
8kbP3qgfT2OjPl28z1qko6pPtRQgUEF0Yu10+07PfgaiLTfCS+N9m+944j4KekLXvU7oOuMhsxzs
X9yLy74isf9ObkfZQz0xtT/rzfcZ9ZIINrMwdvQvNurf9MdF6BwQawQq/Q9MP2pR/60Q+WweeMDF
QNsD8Bli9Dcl35ZalR4RMkIJ2uibad4yBR0Ntad4Y5dWpUlE7+2WdLAzfy/4CKPwStvZBHvDXUqL
Dxs9hVCUHob0xkTbIII3BVmRrY6Roh5AQkTBXEPdT/ACA8DlZJ+Yyi4VwCosA3t5Eex2/eP5U31m
PmsiOfLnC9TrkLM4e1uP/bhZzt0LSeaSQHk0WtiBGfJ9qYzEhXLSvI3ag1Gs499QjCeCW3ldLqjL
kO486Y1/9XHlDO3JLdQiBDEF5pI6fJwZ2FKrKBFEr/SBuCgLP3pj9YIQJ6e39cCoTBd/3rZbddey
XsgCEkwhxwEHNx2wi960wmE4IrHYoRFiKudJrX5n9Z8XY1ZjpZR9pCh/194eD0MkgcKNhNxROr73
kGc/G3527j/pVCTskMrDyn8LKe6i8+/uvf11baOUSXlunCf5+U7FCt2zG3n/KRJjr6J47Ts3sYZL
oXQ65KAPqn8zSczQ14r/Rm5c1FUUby30i4yd8bYEUctzxb8WgLV23ImNXxhszxvf65AfTZlLRqOy
Gr/nYmsicY+S8mJP51gyjJSDdPL9XdKWi/cmhpI30WnGp7bRM2qbSb/hiqzEHLDIAUeD8yQ35lM5
q65RKAP3jV83tTqbucZQ1PHnloOpixE8ymuYGPhMmc1PJhRmOm1g/z5s+El32b+sXTNrJ4yvrcmj
nbWASvtDkBnkVP4+w86c4i643SlxZp+iVgiiSHhxAO06N0qOWtuSEwNW4ECp9ocIHu//tzpwrX46
l2Ow0FWYRzWpxa8DKESYDu0c/S7Cyo4D1QM4uNMsjdsm/VywQsyqNdWmoWezQ/6rEPu+3XYapqy3
f83Hnrxvi/eOp4sC8iR/zvyVy3Gbf3Ytkzm2sNGQBH2tyywEKdR7jMwWXASeDLd1LkHcMFD+qQ20
P0R2ha/8zKANjB/n0PVi8ucvw1T9pnv1tHpNaIRPw/0nOKGPxPmi8nzAnmJSrsC7FlTbTEjBSKiZ
UD/oCyUSQdtie1fM7AvySKR19bteTl86NcdxlGwsCAviltWDvCRe/eyJBtIe3jhMOBkEViiYjsf5
Um65gOQYvB3bjW5tzARpQ33CqIEfyOajeuKwsVq2XwGSLjntixC6d7vhVyeBn1g4jMT+u1xT2ggD
aKituHJdUFS3rE08PEDNy73LzBAyifdypUZKYjP30YYx2sb5uXKgNoAvfBQ7oo0vTuD2QolyrqQQ
h40jT1fVd6/z1USdVFTjsjeGTZoEk+57ANWRaERugW8vIXjNGS/3HYF9m2RGoPqKCM6zy9TJxlt4
SgpT0t3AlYZU1JHwwQIjzYSaCoiAB4nf33mAFcxCspzAmvnOcwwBkN+6eMyrIVmvBnRRYi7TYWKv
icrafq+Po070GzbV/NgQPG4QAnwEDqTt+S0fw0cX4U+Z4tlNVSw0bbD9w1MYMUiNHvu8cfUye6yv
hh2OZlvZHdQyc7szSE50LzoMoa8IlW5/fF+DbWYhoWmjnGG7f+BLAgV2saILje6jq67dbs7OJehu
bsnuek6m0ixpoN1WUZuq3CQBnJh/zb3tb/lbdIAGDyV3M1dpXKkqexAYwLEQ3dAM1Zo271Hu6dQQ
oZPA7Bth5YRwp0KpeuTdUixO4jmVHfJbiqdg/N8c17lvOYccPpfkazTYE0J779RkUf7BCZ2bvvDg
E2FbdeiGhs2kjqo06kP1wkyGrObhK+195H0+Nq7BGhb44H/MICKuOtG/Y4BRv+pmFtyYA0Qq04l7
tE+eWTXFE8WgP5g+M/via65Y+O8ip94iu9XK2j5Xbw0j6QfYzLhQp0bjcbq65Oh0Zr0/rXVcoXlq
niP/cE45CS4iHNuAx59jagLpS671CZbRjfaqdpdcxo41/TncvY+JcqDbKgVTPFlsj9SKpwepsEUB
pYywmYtY+jDSyXJfYEri1lzrdC+zKe3w65TfqknpRO2PgvT1tEE7dNd56kt1hV7lnSxnhQfkB+Rz
5p45BhjRb2LujysrAxuLj3NJWMQALFFUOvNn4WBXRopfzElVetvRIUm8+Yyf8biaXp/HnDGOXvMS
FoGEOSM+l7oERhabOTE/LYZHJuPgLW5CEo+UEglHutZZ+QcvfBYvAReEqIckicw2xTphu6nAzIBG
7n9NDycdiAtBjkx9V8ggZdBQTaVsDfvSKOyYSKpfaSd7v0RHp1yi0hRIvu3y85lca23T30fQ91+f
Aqc+/TNeg4SX8JA4BD/gjANbMaDozOgy+dPS8wF/h3XTnH9CKcJ+uCEseS+sRZ3nQekxFYb993ni
Do3w3roPnoTFIGpiHC4XwQnqrayTbHTc+YbC2E90IX+L7CtSmG+sw+8zeI7Iy9R21rCqam3V1e0Q
baV2eSAFLfYzq4Df30O7YVBDDhZywMz6HizApTZiwV8Lpad1HWXuG9rIMeOJe3C4YynTLb6mUeG1
loLfY9V6FS/PoViEuCy5kwrDYhhmsWIQvNHJ+w6D5MtFGTOgWEen+O2AOn06aYAKIZByL+gXLCaT
kCYjhLsHOVAE9arW9rVreO9iIlxcCGciLMX9eL19PpF4cO0RbkeP9OtujPSZfyiQXMXEdPI51YTt
/Lv8R/l2GJBuvLiEQpaxisyHidOf8l/LV7Y3L4E2i9Hz+ZnHzzE8gP6TcMz6rHNpIzTNx9WJulD9
ctm0PCAQTtH4vPhwomcj8EX9UJNj3JsW+DIFOdnmhuhjCEpIspzcm61t28IApvGyIuas6jf4Pb2H
6r27T9oQSfXdJ1ywV0ZCwM0xKlDYOk/tDM3DS4NhHT2UpTi7RpFAM8+usItSYrM+2asvNJESrv+g
GJPEmHCjNd8vCoyoryxMV7ul0VUXm/YiF9Rs+byjvylifleWyuuETXoxTY/q6+PnDgIVo7iyPfI+
44J1kMz5AmSbqHX7e2AhgnvB6LU4BTpeQV0eIeCGJZ+B2sA93OgHOyDCZ+y03mbJaXpGXRaaqs75
gtVZ0lRo3EkYmbR0XQ8oz7zicbrM/Rc2m7IYgw+knMmpBkTU9z6Y6L9h/ILAv6Z6tcJj2y5wsOBX
F5W//p9PJ+40aBfxFbV0H8TuPrxrQknXD36r0ujXZxF8/JUFPEOr4hTtS6XTEyYYFN01l4TwyjzU
tWv76muBDYtZ6fLk78hZIG5Ay144yjqEq+7xowCDP5ABO1WcvIVYi9pZI/Nu/aNT70yI4/8ZE/Xi
leCbfKDama1hkzT7e7/x9VcDAPft27ywshp1WdRq4PP2x4PIRlIR5PPMux071ke77qslJ94paFjD
8M5+11qAW3UxoCS4HZMl7uMk8Bc0KZXiCEXB5Avuk712z2hPIeJrX0846sSRSuBvzwk1guNQfcw/
hzZUlRtHvkj+FrViDr+HB6rq0jFC/yhTSej56jLX0bEdjaCs+82ieP7JGXrkknIDCMRaAOxX4pEp
d/JlMwfOlQHSSodcmvhObEcXzt6YwN6tLMWODAROIKt2iRVqzvsDlL0u62QNE/1EiVtwH7tzR8yx
+JVtk/A8GM97wBuxkekDUmCDAtQnObe50hw6d+ZrAF1PKLBB4gwP+h4j3G7lOugkD4k82faunzzU
owLOBQbUgDz18q/vJL+OBd5pAwaD4lL1czFwvx7IfjASYwhn7tc08HgLZ4ORWZWha/k4eGy1HNEs
Pit+zKz0CUZjJJI0zYnlsTfcaUtbp9tA6oGFi3rp0lQGFAmGKi8K0FEAyL5NUCCArj9HWcLadezc
ChpNiP5A+90yCq/ZEAlYmv47WHfNXBm859UVWFMSPA+kG/ulMSE+dEIzeNQISxS+Az7nQmc3u3at
nraEoSaGMurPSqKvUhz1OiYhtH+U9/1kduedHEfWkjjV9O1skrecAObMvL5VSQY17Bo0SXqODX5S
w8pij+hIf6BDAxQzAlMjm2bYJm+O9LwADIILb4/ZjUczcJ5fL5056azKD8PsyT5bFssnbcCWnlcY
6LLkItry7bnhEmKR9GMvXUeWsk3papnElRzW3hLPI7ztjRCOZ5Cd7vYZ/Qj/prccqb+dIDLVZm3h
TmC45Z8jA2GL8xOHk9vH2skDgCphw3CMsAOsxae9Q5nNjHBXQPLp6/B2VusbHjymHI1sZvR6Sz6T
nVY6Wxd/xJKrdYmDdbLOgbfmZrsRHljgtuCMIHeo8VPh15MvJ48ixfEGow156OGg7BHvMQPdGw8v
7kvnn0Bk+SAgd74Zc15W88WnQ/aC1vhLUITkqOsECO8R5G5J9rvEQ1BggOGYnVMry2qetvZ2xYtw
/N31V6af9qbcMP51Vn4XiI7+VjrdcAh3P5TUEBf4CLHyJHr/QNcVyAWmpEVn7FUtDCMfGfQ5Y0lk
DevDlhqwOCXqV61Jdmb8UjI/g8L79982JHTNluOYKaazE4TCLNXZfjdoISd/XJfDNpvblIw38bDa
C7GGpiiMkxlEgZHqWbczaYQ+FbggOQcbNdUToXLYi/pr/PXHgAr9Gr28hmKdZPpi037YRyOKJ+lt
c3cFGwRDo3fRj1PE63xXj0SYxgL2R+jOmy7Hxe8s+1lQJXWKwAHdp4QV+o2wVyxFNGTwKAtoCWZd
zNXjvq/qWo8qpQseE8Rtu+6936X/DCkKzr+Emks4TJoLS+Bh8jwoWScK8ZkiwjlNNz75iNOBtTQZ
clpvTdQGcpKRynpiuNTghjFpTdG67Z731HQwvUMCyOxyfJ7b3lRccXmWWcsRMqn06Wb9c6GWLDoH
yVC/vwksDvn38T6Se+a3K9QcZHash9JaY7DtKsnqjFWn7m1SBs2l9daGmg6lnMKegWq/K6ZXihjm
KWZFsvqbQNmBJUnGciXcmzGYiYkRLbIUNREiUqr32kb5GUGNxHgX1CdPI/Qi60z90mAmEUNfghvS
tqtrXJAetMT0qvFVVvyyeTj62+T/3zzJGcT3fFmgjIdeICudzLmyj+RrVa/lnp1noYm89IipnAdH
bvJq2KSKVCxfNZ4S0RfNXyzEFq5UagQ+W5MOSsjA8mPS3eqlaWEXGBbBTYtuIxaEP740bWWPXtF4
gO17hXQSpg7NvNrSIt3o6Ca6UGyowOAyhUGXFFlIF+dH4rGGdZtS5z9V4+MiA5k+KEcr6x49QcIv
nuXxOE4tLGwHMSYMyNY+dMctPIWzwi9hsYWaA8KoCVrQ/yY0SIIPm5HIxI/MgBf6Tyc5IruiSyI1
pTTJ40L7ndvTCemokRTZ+ZlzktIV2VFNT+q3sW1WAMPgzl7eS0zR+6aG2hZ70haRhW7j68xtl4pf
dPts2p74F2ifBUFQYg3jmeNWRXU7yAtWTFo8a7T6UgANuurHoovfOlsp6hrIMNW9s+sZ0WGKnkw1
O/CtYfKn+4e6Gy4Mps9NEXYRuB7mNXFETwNMgIzktRiBYUETI6IdDLLDPkUlK7ky0oJHP1TQAssT
cLXsoCjIJyvvzEBXk7F6qCdQRETu/ay87uXdowurg8bIh3mOt5KWPULT4Lti6IqTTYIBbZ/pU3XL
KbsO13N//kXEOUayFOOnO/0pkmn2/jZaTIuATuC6WjYLRiPZ6hsZT99lEF2bl25RL6RYkDHSBzZG
R2Qyy5azoeFIak6dpccAWll5Hu1APwasiSBRZ5Z2gEtPfK6S41gY8zyBOhF31uAXJGK7Ger/enKn
koAiFGdhleDr/pwBhnSgNBP+VGkHaNPbZswe/UUszbuEzWzo3+hyZ5CXtzlRvM8IiPpafrzkk+R6
cfbG9FHt0Nlbj0/djZdxL3f7jvtg889xgX0WYzjT+8vDDFqso4ywTOgOubTi7VjO3vWSeHhUMp8m
gKxjIJfDpePsfmrn9VUECn2J1SJBHZp1PwS9s1Z8qhUPyhhyEtZT8p8ajSrOIf5VLSPInqYJNxFc
wkHw/uIcN7F6Cy8JTBR4fl22ZmFVtezugccZPO5LF92TwK1X748XnVomHjbTBNFpOO+qX5qTHZzv
NK8FFCoErBO63wF4oRoItq+XqGPxeD3rknrTydkBOyixboQcgb79ux4hKoF5u5HN8OcCh0HEDjV5
32dHdDi3bKtndoVFZsD3qoDphmPQBMEQt8Ks9nRSOqQGs6eRN+df3h44TAYu2IJSlKw7dGDpXRxt
1YsGB3WOWETMn4DsGK1bEC69KZNE8g4KSBE67zgMaIqzyQ891BKFBJCxexPYBzy0mbWAKNjlLlXb
1og=
`pragma protect end_protected
