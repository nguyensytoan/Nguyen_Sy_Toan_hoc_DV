// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:32:01 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nCSS0MOCAk4Ux5mshfsC7y+sXDQhObKnSTVOXiY6j8qjcEwSiaxQoG50eSnQf5VV
/fBiFZCyP347bP0B4nfnVD5171Gkfq3+ta2dIzRKYMT/uNzEv5dR58Iq+jM5acRK
YLBoZl05/DlJ6mSUoeDETj7FtZIfK6HXa7mWoUIpLGQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12432)
b5Gl0ApK15dvXKhAZP5e/Vcrra8kNZJLTuRAHWSAXFxckAQwHyDXxZW15nbp5u8/
KKWKcczEIubcdi2gcd+kmhLt1CITI0/75rDOwHP4gsxh+0Aw/6SoeSeYxK4CLl7n
7r1/PAPcrqEkANcuk5qcybtOMgX+1oXstET24+o9NLFHcPVU1lBYJzfsApk/TYsY
/dCCh2pCgnQ1UYjs/MybisTV7oOJpoE0ZPTY6wFdXcM8y+mbfStGgRTqAR4ERiqz
eOmm/U+MpofEPvwKjXM5KTqax8sm5SbdWYfxoGUWDfWGglGXg8/isp7ADRxHJhWU
8CpWrvb9fGGoZ82k1ajRewLH/+Hvc0o7yxY0OpNnAOLj3920zRtgY7YJNnpSHB6I
hTUdgIRGkylGmYmc75U1k0c46beP0p/movAABu40eT3gc9MXTxNoGg7OaEVVYWr9
iQlmhh2qgL13dPG3OCBxzgFrv6H2ZUURp2p5j+GprTbvVNKs3XgjpXmA78X0VkP0
HG+giRDYC6dvhOcLzkxqPmlNN9sYyJThjfoBuv2P+DfbYw1PxR/9qKugCJ5nIO6u
hOV7FlcOcZq5uvnOpckbqsTwACbH1oDcEEWAhTrn2wun+xyFvcJwUIAeGU/db1j7
pdWpvcrCvhqdnXevb4M1SueaDOJuqXXdCchIDZ0/+qQfCfg6tOvsZZYraHYsVOZb
kMcDYThUtiXys3lswnGeGYuW/YF3wMK/gYcuiAZJGm1/9QE+jp3yG6GWLH6IDhr1
Uo5rOwOlMoi+ToyMnSDZQDq8fY2vWC4mO62gS7tlTkZmfGaTnNfnKl6xMwdBFtRD
TzRS+p4Hxb/bB/2pQs4BGysE9FX6wFuU2N+5WAB0LB1oVb2iJP/Q2RiEMGOY/Lh3
Or4ByZwqVA000SsGHskJu7uo/5ZISRrxiGjKiK0iiR49sPqxLcAwzv4Mlsi5xNwu
bMGkeo+45POSku8sG/3VOCalYcMj7Xp/4on1MfF7hJ9SbZpfOmf6AhJ99VldHMnx
a2znMUzE+H8Ns3VmYQv2tTyhwnb83eW37Nvt/KQ+wKHrpK4V8t4SNGI9PnxERzSG
Tg+E0ao1JbjYq93HialO9LJRFDp8ir076NGLIxPET5k8ZdTHnI0TKwvCzPOirw9Y
VyELsIfL72CZGSNu4182lZJTSHDixFultfUURj+eQvmXNdt59La6RJ6+4qRSYrzQ
BrprnpcIhwP4G5rzAEEC+6UL4RR0wjetzriRmV2jUIIZLV3gjl/eX7RkQdYlWIEV
1H9DC30p4as2bOgkRFiF7QYdJD+eS0MUsqPx+Ueq7CpAJuxCAbDnh1K8xgqor7kw
/MO37jazcml02e5QSTn436KNhiatbpEP9vnmPtJjzT9mnPemsj7UbtAYdHrSU2iv
eofSg0iDWdydU/82qVovYk72ahoJEweoPe0xIGtvEKeAfkOddlutJ9avOo2NHPKQ
cdWhb7MDs/v0Fr3+K9dAcq0SFNQHOjinLyWIIw3bdjhPjgQc+vKj0VV/QUtw7ucV
Rh48ppj0e58HPt6OaRZ96lCY/3s9dbJzYl+LSaq51doClwg9lPgVyNVDLPW3eJpE
Q5rUCXOYcsdpFGLHqCjQBJa/ikRGiaCaPbA6YCLQIpsQUKVqAEXidN24ZYq6aD3/
uCMys19ZAatV1KAYYnAsuInyxIDeNfsJ0y81E5P0fE91R5a1RM1WZ1mtkB7hMUSY
tgrTF1Vot+i2gDx2xI3LxyyILUPBTpSV/0nnFrA1KVrFNjcmqC3Of57AiT9/jfMR
cu6QYe/h5lJuSaCrQMb5cZrbDxjZ3PfwEI5HSPpD1vbcc61cdzikPg38dsqS7pGW
BjtWpz7/hEIaPWIQDpGYLoId7pmMs9etYD0SmCDLKeufzLC38vPcnWd7RGjI0OvH
l89b6GNPjZCrrkOgzwnDgghcCOLJ+q+PtAXyvvN8qTcfG+qrtmgbo8Inir9QqyXc
5hgjl/gYG7uUt1hu+X1P9UyYRhMSDMrNyp35jA8EcZfq1GIO2I1+1yb16A5tptbg
PkBDwRK9NR/PAi2VPX6Vf8s2/7j7rc6XR1dHWnriJTnBLhC5GifbglEFieW93gdP
kbeixtN4m8cSc2G2OqHxdBRE/4UEozU9QVpk6/dxkBKmShW/hcTy4kux3MhJgkB2
8odLgndhwrqgm2kNt7rx78XXrr6tXoHYdy9HH1lk4rLOBqLRKGUiJUFCGYH6q4uZ
rZJ7Pmu2PXmQpK135DG1fhFyPG1TfIBeDymun22EG6GCzrCqJcv9/kZSMEuznu44
ttbUO/QdlbfQZch778JMFAot/JsmRs6goIDIH0S48feu2FJuCAO+RdnvmSZ4yrMY
7ZRXlh2WpeZgEBf5gt3/mTHcp1xJOnhIAUeRGDKsutiJFpODfi9hRV5ksuho2+Mi
uO1tal5mkjb9On2SSnaxki3R41zhC+sPdMVTQrOK973ttGoxx7rPXEh5iWNUcvG7
KzanglSpLMOOu2E2ppQleyTnyv2WWExt1numraLhldopkwL891u5PO2kWjKxV0YC
5kPGlUfnx9gxaxhcnrslseXr+Ccvu1fVwvLYPHt6sI+UV1f0e6vM6Au6dzcibxCV
MmH4YDveAx3KuYiOYV0A8iJZ9Mr7zVgztyqZ0BmjjRRvjPB7hsnDI2lQ4gTbIFxd
Dy4JVT97SgXeKrcYo9/kkY0mh62dSDjUj/dE2A+Y7Pvid9beaGnKAYpxJX4sC+X3
DWBnltTdbrPvshGYHGOpKzojBcXnlCZ8JE3dl3HHTy9emI7Vwllz797OaYjxkEVT
5CJxaM1ValOX69jy2anYTjqjHxhXtsYnQ6701qBmlQKNi4IOXrirMMAkCzpgBih5
P+b8DLdny3Z5JvxiEv7ljSVeIxq+T/nzeb7PsijjVfoqB44YZZ/NXrlqomJ4Wbho
0sFCFCFiNuAO8bOrHuLI2KLLOGSGHk3Bj8LyH54J1xbkmoXXYqJOceIBDpvVxqJg
+8Rgo0kWvpWNVcMmOM+6PWpApgVZZuEmxhWdJVwT9ecTM9ICozjJ+ZtEPfN6cRc0
bpJJ/quJWwvllQW8ul94gYGtSu8AGUoGbXSj8YAu63BBhOUrbuYXzHDw9jddi03C
hoIul2F2ufszXTEXUDICfOlQ4CgadkZMRfs4KjmsjpPxTsbCcvDo+6dOY4V+kunJ
4Wvmtrx+Gau3/n7sgCZWjofDHwOytFhg2i0FC/z2xav+44BctFIVt4jkNCcDra6J
qDaT3QZLfaQqNiXoauCTWRLwpTnc/aLhYTJpOqTxcvbsHUK1Xhpxffam9Nup6wfh
CmIR4yF9peu4oUYxaFXNRG0XquuV9RkP7jTxCpV97aIFF24jJ+OS1ykXIqkVDnJs
LAJj3unLfHRECAWOSAk3vpqRw9G5J5jqZA8nf+4k5pXW2DY7vjEgJjokpn7eigit
a95wpgM+NbSNMztVpuU+AZjX4ircMpW2N8LAXvSIa1sxL0WkegYwyiD+wr7IE22S
kZ2yZWxKRmaqiFlGM1HzXhzw5qd/rzfIlWhn3G/dzTT0WKS9KcUU0eNRyfDUOlX/
aNJNmrIVtJjxMm+0neLS1n5Ein9whKAAPTH+Aa5fIa/7yykVFsCS84N8Kzp3Z8uU
qjG3MVFpjaPAcoK4+JFIBIaFXuHoZNXPUik9vSQOrw4Qj5S4+D8QWub/tU8zT9Pq
b4xdzfa2Jov/B+g5gXYbqlQIibLmpYye2NpNZV4NMrh9miAJT/Yrpm98lnjBTdMb
TqWWTtC9KUGNKYm4RvAKCQ10UyQ5nLYLiXKt6WBIfWJ8fM3O5DSc0h5ZzcwdcIGr
0FH05jtlrk9f7vOuovu2KCaOhOi2AiFHWeySz1TpruFe9eHmXuYpwK5rUWSCrZ2a
Cpw/rbdPTHrQHXJhs4NeortGZIFC7TNqPC5GZyxU3wtDJQy/d5uhNn3AIbvJjtZa
ZfRftWLk8HbiGAEKj9hOSBY15kWAJlzl21DCuYshmISIJsaeuR6aAZeqUr84nYTK
zyT3bqLhFa9kCc3yGFD7ZgkX8CRUr08TczkkDw6ZgjRBhoFxvlyJzMHhZ0jPM3XP
x03mcmmOCL2tXPpIOd/SUdwuB7bwPlSNLmD3RazBqE5cNU0buBeTkO0d/E7fSBOb
1JZDM5varS6idyc+w8XgEOJJ4HPajbvHDzGv58bUih4QDjjCWnYNJdP2zpq1KN9M
PGRVEqBcRU5YEu8a5q72A96qf9DThfqDSd0Gf5lIROThaeh24JweQp/u4tt8TEBy
n0Mrg2HWhSCzUqUJH42YsIR3HwmtrBXo7cIGzehZJ7lSq6su/9bxKtxh5fV1Tu6G
NPhDa3NwoCtwQ+DHoSPIsxUndgzHG+OIqtIzaRBKTDig+jP/PASRaiDyqfSUOhDH
CU0yoinxX6PfzsJHo6owxoF5Y4wN4HuzoSI8D2GOjUqGhmsa6jNaKPBRjARYccxv
VuKDiQo9N99faxPh0lK8JgfrwhrOhfbzgpa/ghBduDXTBLQdVSOZfFMKDpj6G5es
Af6IulBLKgVXzudydaZmxsRI2z+AzJU5pphGgWaZGxoUdsZYJq6nqKmINrMvOExL
E9NPy/EO3QWRLET28vdD73Mic7RR7/oOubL+BQ+7apO5vQian+I0i5q4H0q4WarU
7o00TtAau/YOgd9xg4ktO5l4fmG3lGn3g6/e3dns28WZSoIel6Ub9MY0JM/5FOtE
MEhg7ET2w89/caCARyvlON0oPB/F/FY3cqA6ZNAzQSI9xdkAemAI89my3qmazA5g
baKmAkMKdgPhLnIWshxZXsPhfK8xiN9WwwP/MvVrhPnBAGmDqfAsgT+OFdbAhFUK
OCeTAuPbyOjXaEsOGeUs2+FOvY0HDmIakwGohC1+MU08YQtrDM35P6VTuGCTTz4i
Y4QwOXKs/2KyAl9u07X9zpWbeTYGOeTtbntsF2Kb4f8UrDXnY//kZxcDhTagtM9x
47b1YOngyPucaL9lDEoOT/jZTuz1sv50E/38wNMmDDuSWtNUAW3vqEKW04e/0cZ0
tB5pAYbgzUP2W2vLUx5CDz7iTWafgjpTmLxzkYdq8goy6Vto03PGGtam4xjGFUak
C0wcJadMlnUJKNhNYdsR6q6yLhVr6OXdPm8NDxI9nLAOaYI1yJ0IBLU6UqeQ/RZB
1nuwdWoHuPm+anf7Z5geYtXvwF72lTeXxbGBk+XMeBUWEoEQJbgBCcH4WoowGPOk
bQi/XeWyY0J9TtytnnrA9CDOVOFITdBGLuKAwSFQaXjsooX/0sI7QLvN14l1QLYx
nfEROS+CSiYWgTHlzBc+ignwnYFLap9vOZsZviK/GTjQ3bRzg9hhN78muBrTrslV
pNbV+8Bv8fBNk6AK9A7b355Y7nEai4Yt6DpFs0H+u4c/LBcuDe098YJ6jezst3bd
qqGhWPKF0v9S8Wg3XzIqBeNiptfO3O8Fg/sSHh2nVjF8iY7Y/7Mp+InBNARnZCTY
ezG4Ykj6E2XaPTRrvMaiXszmIv+cITlLe77uX33dKm6CX3W2TkZdc88NdNGVxXRE
0feMSq4670wBXMCSjkkZditc/Qw25ufo8rdUJfRLePA8AP0UwYGza2SQgeqaUCX5
d3AEiVH7cHv0PuYcko75O2flknOgwwC8oxUZAmB7Y+ymKpVqtFqyALBYNYCVnn9W
nD3I/+XS2ShZeAFiRBnE9X2FueX7FWc5uJYjKPnVlOdmwDOwuBoe2M2I0X1SsCot
q1MIiQ2aiHgcPcHgVI5rlzTdDBZL/o5IiHn+L2ok5NBKYpxNHvNpF2dHfHg1tx2Z
Tuo9gEydLfOPBe8C93v1kZMTgn3ToDy58cLI4LMXOuZISX7CSOL97efEyjH/QLKx
vVyWrAZ3v5cb9hh+xSD/HASo4BiexwYRTyARZYpYt3ItfylUx1n6pLWsdKewLlhJ
2WuTI/Obn4qgkmjtjVUzUpb1g2kmbHmz0G+skWIc0hhxiAd6tZsoV9AbvcSh8CWD
A7rXk56gG7U+h5EVquGp8GOGNnCO8UtmG4NIcxJ2bK08FvTVhh6RbDLJ8HBidu5i
vzAcaM0Q+ODuvYf8LOThTbRRAcEfbli/IysaOGNjKRNt6xvoGK2+wIDLncYj+47a
YlMdtg1Gk+Ng5+ducFBL6CENX1e2FZN9rBKYVb+WaJ5yVHxiuP/BbgEfBGbqfFJT
6iMJbOwjhDoEUBtcem69J52Aekq6UirLdxplTxBZixJQeFNw/VGLuINto3Gc6etb
W0CsNVKg2AhICuikQQVcs3eZA+iRkatRlmEKfq2wUnenHEfZgUxr0iB3v5k6wnHt
FOqhlBgYPJQFO67jJlbumsOjaE8OPOtLHwmcePJBxStQxLDoKJEcBbcfDOsk6CQl
tPyX2w1RlZHtRlEemqC025delzwXT3Vf6nbQUrECVUYtCoyaUihWWQ9zyWfe/wvJ
1NWiLrm2r4QgSYvo2GGMSGDZSMe4AMdn4ZiLUXYqh5L9pzscjX3ydEJtiKGSKcni
+IPhS32tKEi/5QisJKlcv6XWaphR7CaT23qjCgXsUS6BJuGSP9gSmOX8/U2sNicl
7OKSa+nc66eHi2+ZuXWqbaqXl0gdolsIeGSZDSMNVrQMqVdUafCdAQ3JpHsDcy1s
lv7V2GrKUMvOXp40Ndb6RxyUW9502BtelyiJEr5ciokZ43Z5wLiQzpdQLetgZHjB
92GawO08U8nh6kk72Tj22SMXFkMm2mkDZdOadopdOS+J2AcHjcadLuJtZtT1jmR8
FIxmABC7CK4djzLP3KR6Kxrmv841rkOO4Tnd5ktZowjlEZV8GWJyaTJG62oyhw9X
ztdTIdc5uL79DUmcAL6nRtf0oBySZ4qqgcZVGdsvMftqMjs2FVutXHTJahpT21ll
HhSEWfo5Fv02QxGiMqhzzPaG3pHnTKwCySpWf6QhtxqN0cnwP8Hj8e7bA12n+/tW
QQHVLgS7Q0dnVYT9JTreFB8KT5QTeKhl/LNqhpTSi/sgw8rMYDzNLVo135OmHDN1
IjuPSevIAq+nsN8f2zAx0nvp2fsX+lAmkv1y+R666OGQe0zhpkfIcwUQtUR1apx3
509nybO2E3IChv/HyZ7pLDREYDDFkqmI+brxqQ5czZlR81AclYBR8TY8oFzeWQTH
tCBbhcgURYnKQkmX2la/5yfy+aRBl1b6OzXWH9xln6NNdva9dknjVUoOflnuDU1D
dyN88UPFwCE6tihgWTA7nCljV0VUP/BUpOKunNRGYyN7T0fd5HI78lDO/pNJpalF
oAB7Bm/OPBjsVJEYMLhFZVjNAUjZ6DGhg+bf9wxjZJTANjecC3vNpGjwcDjfiYzY
RxQVvXaVGuS7HkdMY/U2kjTQxJM6SHunQD1hqSJbgDT4W/nFmeo6LWndbg/3uUuP
pHVYeIfn5SK8DN9B7xe6ES3Y4i5nhhjq84+VyKlL6t2jMty8gNzXQuDjr94j+VCQ
WtEQ8uqLzRVuWXnLEaUlaqXAMuKFpIV2x3ZDykzr26ulNNzqK422wiYcn61pjLgn
HVL30bRMxV/Rg/U37LDNQhFKoARPtTOjJaRdnWVz7SGWxZzcs/w+qgpkc3I12i7o
K/w/2Q3TULUAfwAA8YIHpBX4FH375npqZz4BNSBW0daEEpLfQWMHsQz41y3+mlh2
WyoUhUNSle5kL3+9wTDT1G6GrYUkszQyFHL4XBVaC7BEaGNAEswa7H00zmnV98G0
RGn2el9XENk8Ax/Dkm5Y0kRspMV4eVyvofup/rSVE0gk5AAethYI1VLgFgh+t307
4Zddge8H4PUR2IZaHsQnUjkjMO4yLmSY4kGazJSmLqFlfcSFYlKRG8lmJjKPYfv4
vkG633xSszfwvOCm4LE6ECHronFGlKL5FIP/reUgNnwbqdpDrDInytcv+Vyr0tb4
jfH8Iz7VXOfUJeKBTcH4brzAVbroOUB0mH8Z3oXxj09I4vTjkl7keGLcbnBTHbA8
5mhP3faIA8MYHxyT4mYOJuGXRRTpNFqYX68VvNfbsclmdbFlkPzZF/zc2Zap/X8r
EoPmqa8LREsnqtnhpvpdS9hFBoisZM0XXCeIe7kzC9PONr+t7j2Eel+D0lYsMpCH
4I31rYAiBIUPzFrnakCX/ISisQym+QpzvD70FSbfHTepj8FaLUiSGVdGvtImwMKz
RdQLTeOgmGXRzfvwRcdihbyb7zJfDE+29DPqQ1xWGm8oej0N+McY8+JpclW/nU6R
fn0ima/YiOcDRlvvuOENYi4+juhza6Gb1bOw2CeDhcshER7bQ79SLFpVnySmPIWK
b9niZPRRUfkIY4UME5A7RG6GwXjr22+Q1y0AOAYOTVvIV36fR+zgkvSw+wrO7SZ+
BsI/TSQlUOUvI7Qrkyr20f4CveS5ytz1Tw2XFpG2hmd5HK/8sQo79jaN9+wZib5x
E1ypIUVOoy//DcsymE+TklRbeLrzGA7+1z3tGCs9YwlPDDuk/XkFYO92+hFVBctA
wykriAaVFqJENQqIdMEeU6ZbaQ8bHNTNjJLV+x6isegbHEwV6+C2X7qni8pLB8fz
qoGrtGIsJMm6vjpiQuakvADCgJeECmIh1uTblpAwR8HUmpfmOg/8WtaSNqlFqCpx
0ZeTvzYvWK5Zwxwc1TQlkxPXeXXHw1lew6hExbLUFxO46pxDI+Bo3MiKXDM96Dqi
4krEL3i1RfZlnkXEBDCAaOBIHaX+ObJRA6+JsQsowsRbW6ie9qUbYLWi2mui4g2h
svGrQpHJ0EeALFnzADnypQ2c/TUODDK5uYHQltGzMfL8/k/J18g6WIVbp9mYuWaZ
CZc5jrDVgci2vib2owmTVhKufl2AW0bQJIAv/fYRr2Qheiyu3ixcU+XhVzOjAx/X
QG0TsZy8Zp9Maf7KgQEACGTfO+z1SKuBDynrOQIbFyjjkJNiogl91cHD+wFWTA1v
xu7I3lixIRBy1IVnjNTZGzkUie2yDOrJYQUDJm/enqu9xFxxYJmqC0YB1esN9eB7
z3IN/lAeIgpK3cytCSZVJaGB9KcXYDcBp6wZLfzzBmpq+DmrlL9rxvAY8LbSw+Wi
/23A6USW2BNiHIGSm5uSXQ24vTs0l8byxIzLpJy+t+ap8HSnhEVXNSVJjrO7zQxH
OoVPOQhwhuvQe7PCtXywBeclcBdSMZqhntqPPx5rx6709ahgXaoSoM6TPrZh2ufu
9RoedctXJWGGJAuKjCHWZkDUifrHmZMWaQBbgTuPVBvMVJ3zLVnUC1hbD9AZ2O7h
n8KipyAxQZLSlIjzYev8bqaujxjho9RAlkQnpJtGwRbsvyqRSH3/dWFaSpUnRsHg
VwOd4X0iHbFZfvtvBot9haf9YQMHC3ABtmhKgyKEc/mUNsuMHuJiIy05VuzF1oNR
YgS3O/MVguwjatZHBe+vsUV9A5DwMDYJMsb4XlgSYMpLf49vHGaKOa+frfGc9GBP
1XLnUWMJgJmLfO9nECWaITqDWnAWhqpW1C6nrz89r+WnFLeQzb6Q5YoP0hYj+rE0
Nc9A+fqmkXJmdHrJdkSnkpjXuBdXkRf0t9IAN/v2G4GVlNSrUUBJzl4aMEn6M90A
8m2bzKb6SA1OF8pSIuZpzKodEf2MccwTsbPedMA+lKbYIi85Pl8WuhAyR24ow9X8
1RIT00d8A/CNLaT3rJyk4ewnFabFO3S+cLUgNEBFBKKcZqIBcgI0k6FZpVDZjBbO
C4Aj2O5HE8cUe01y2//4brNj8z9hF1XOUodrVEGqINcOeenvUcQUlHBDEBqrdJ1t
93j0luMLt+El8ESUWl1FN4AhKjK04Kflh2b7tqlCkVieaEB4z1l4cnUBJPvxhRsU
XpujvCB08sUrPblLeu8Esrw7va2j4XomFvkWe8MR4ZV2ROCgAo145sHbppsV4YhY
kt7NrdufT12FBP3cUCH7sBjSF7ieaG2ZGqgVinkeyGckGycWALNsfroZBN/hc1LT
vXHMPFctiBvwb8R7Qh3/YoniRkSEJzyd7DDu1ax9/pKBLQOLiHVJZ5Vle7hU0Gce
EAAZ1FWbCjB4iOwSSFO2/WtVKhMfbFpz4PPRoDlMRNE5HDMBCW3qbw6vPuCnMLKG
E15JxTw2TIViUdSFPQNqiu12BnMsLtC6wF1Jr4swf2Vb4wBnUpkI8M3bsNS+6pxu
Rb7QKhkSRvGYdsHXPoYTzYl1XBHanW+5ppv2wzlMqdGFVeQ8OxDGO+aKM3odvbdo
Z07VqPbd/kI5ZATOGGlmt9FVoEidIjuI448F1AaYVe9bxA1xqjj8oZj5Gb90n9eo
+JxY2RAzXFUx3O76v4OzDavE2CwQgOQ/b53JVNkZIOBk4ppGW1GhjmeOxINwnili
9WQUywlV3MLVn4e9n4arbjuo5eHJG6MdtzmcAf/HflT/LFwhYcnfx2OHQmYkg2DS
jaHsDOZWr668CPf0XmnU0UnDm0A0mn5c/Q8Vj2FkLR7Zg6ONJjUF6Ak3WI0CVqvZ
kjby55J6LsCdcnIBUXFnJG18DBIAK+v5Q1BGaywFWPWBPr/sJMU+SccpUOpSNs+t
IuZQwT0AEB3hivNhZpdIIfFm/gf7RFGz/TtvBWk1O/0v13oPlT4fFw/yHBBnJTyA
hv0+N7R5Qqi+5lnMLSCCCorgmmyUPWVKSReHrnPJOuHb6cvGYnnjo3QoAoVT23Uo
8coSUrirdTYTW2WE9BYVkiAuf8xf5moYN4VnBBVQdXrvXViAftuvnnr8VU+wkkNZ
6sESHlmOCpZ126D6WgT/roRwp6aduChHlTyUnyX/jBlu9gD/aK7/V+8l57qOehcN
jiuYVQhJvzzKioVj0dyZg8QEW89T1G7fdv3a4rfTMC5k8rMmVo+925nV6oClvMqr
MplHGNO9r7b2o4K6IT+Gnc8af2Ygxdpr6ZubG1ix9/YHRppDG/ZhGKjq0mqA1ti8
R86U3aobrH4n1drPEx1fTWRrHzsjCrLu45+R+4YRWSwswm5xRha0+SUrDxqmFYwN
+OGtZO4tHJgqPgYebyXCVw0sxYaLbXFoIQs/4tIpfKuKs4EbVOIQmnBiqquZFzTZ
WK+eE45hbQmSmqO/XlagPLgh6yu00grRwNfQ0KNo/zPwSce4E0ZXAPCOMcpATEBL
HGeCwCM5QVqqOcSArVkxFRpCAvABhKaExOpTct3MiFUWIe8IE4lTaSBxtxmagM33
mkXmtzNqDqjP3Oenfz8ByPNt3et7LS+QgxqjJeYMmSrQYfEoK311jB0UcTEZEJCi
WaW/HFRgQaZx+zgo0NS5POn5JGT6VoKt58qV7kQ9ucz39q9YIfXNOIaUZ/Rg586q
aHW1kSno/YPyYnQJC+zK0G+sA1Njiyrq3rfMugLBYpom1HdwYuf5Vr79fLT4wSjX
IZnBiyDYKCUMOY9vyjquCcOMEnzh1SevA7PytR955uXS6NLb272k3BsXqUTfYpJ6
9PMQ9se3PNhtLgWaOkc/0cTl6hKVq88s31YvnxqyWF0nLi8LpnjN/+7qbliWrtiy
mxHxpP11zOmmu47cPVPCuAXvKP/eX+ASDG4gkt8H8PQSBbhlk0D5sZPCu2n3GgWb
TV0/CGvX06kkqNdvy8vff99gGUphbAg+o2MyMx1nC+9dJCbcDK586iNKGwTaTFEl
YvFXo9chAePihe6Mf/1SCJVHZSJXcaTa9D2h1xxosVLPsB2NDPNrt+G2mgqswuKt
+0k7OXWEO2UII+DXwAOE7IeZ0hGbSDc1vPAS4HGjxapWkOHtK52wv9JlPb3pv8/Z
cilTxR6wxAYFXNyiokFfC2486CfUgsEB8taVOh/pd3J7cm4KOzei0mTtGK5WQOxw
TDgY6gECsmVaddR5CI5vl7gPrlu46Is4cFDt74gbzI+2PtftXKroN4/EQZp/Sxcj
8upt6u8Iwttod26Mh2R6LfcFdfdGmZCHI24NsngUZpRs3h5fpQuJ95gIuWC2kohV
U5M6oR//arHZK0pfDIa9OSOWqKroXXxeKuKvSHJ0QQ1X4+Fb95DlHwGBpXT5YT+T
NowPWupu9c3hH03we1FqvLB+Y3Tuwr2v6A+fyVEKj+pNAybXODQvJXds+m2L+RUq
6tHgoelURsjqDOYsjmEa+WXTG3xmnqKHorBPJ7wB24ru21qvFQIApNvzVCVo4Ix0
Bgdc2PtU7QwVcChsZmaA2LDhbVQeI2H3mhnpkCBFOxQOc/iQgXZGjVxwJf2+Sf4D
y1I4LGvGLQPlWdXgSLkI25zTPsIsUNp03HtvVXHTkGU7qeriCDqyvHmSnSh4Piuo
3fKU4T4gIct9qkbHg/MuNguT1c4/E728Ivu7cXCcyIepLXQbD5Wg9Rvlq3w5nvBc
ObnmwNpYKVZKQmy4Y5GOVuP4KY7CPcnVCUZSBE5tUKu7Y5jdF+G+jdOoHk0M12f2
5+2pVBas6SGl4XpeGktdqbrZIHcdqSWl6MkM4xTEZ76G0TdZeIbFpzHcRGNto62y
5qRSqqsweOiLj0vzMqUa5dvpOZQd8PMUNlpUHW8KWuAux9vzXKtaIR0/c18fcAXj
YspQR4gk/hJ9IMZLtrzjJdu6EqUgjudNroJq34RV0FX5V8EiIYufOTrUL2ZtSN5E
s2ZBsbonqs6vwxO3z9/GomKFOHPv4YApN/ImbGHyKieAvsrd/Bs8RbIE3/2u78Hj
QhXNCgLSlR2pizZwxEIVRUfBlNRMbUe4QwtuNOr4iOWYgucst5PPyWMaNe1kdcHZ
XTw2BkbsTPV0DBEaLrt+BGk67LjScCHenSVwDt0dpB87zikvJLjfFWiIOsh/nzua
DBFv3iSLIQby3WZMh4w4zo8JHAF4rmEgFqUzRZdb7whxTh6s6Cs4bzFPsvztVoay
3hcUD+fa/ToEADdUCXBQZA65XcMzHcTFCJcxHug0tLPIPGF+IIChdS/MGksNaLg2
2DCtxowIQZ+3UVGdD8gyNi/ZKMNdKRXuY+kDl/0VSR0v3VxGSP9/tPD9Ex1ZBwoE
MkzT+4GT9tbrpTIocwFAYd4GTW8suT3hvLZD/SL+Zwd9rUV8xDKm8b6eFaVrH9Mp
1Xzcx5xS8QBHeecfL0guzKQWeUgj0EADcY9RV0d1+RgflDRcpaRGXVuE/j5EOyHd
fNyp+jxqLOnsgF+WaG7cerZQhTJ3Pk20WHLWqmUVe/dwRJ1gYj+a3Wq3PbC7KINV
dFUOA4ufIGGmIyYvhCLlglcWj5N6zPoq28gHm6R98cpd2nAm9RBZ6QLl0+l4e8/e
8iv7lGilu2HJ52lmDyaYyAoDweYz6aFhHWbt/GsPLFuASh3P5ssaws8jkTUijV4J
fZJipsJFf23smYEhvMI/tluGA3Tx2d5Jd6uHMTwWc/7X74uiuGrVDDmY1N4Ig6dR
KDyI6ns7LXDxyFSo38Zd2j6EX8azxvkK/sQF8akwDZO6LzZmgEKYp0F3tjDJkCEj
C67M4zt8Kx14ROBzPq3tYkih+KbCG8z1rw9PnZb5SLc0jeWcutvhdOmNVx0mcEAh
/s+OgC4bczzPfR9WAjqDZEUzcOjwOPmXSZsrfXB+3peRHR11Rn6BwExYoun6AYAi
8cVDcklaTrByWxlvdTo50QVDiLCUpeFWdNO6meByujnuL8TnA/Xaha+GnGZhh7BS
Z+7MVJDRj86UEX0nM58Tzp/CgFY5exy1bjhWvn1eNeHTczFzDF9EoDJeGHUt2T6N
wMlRfPwmIN0u7SXkEVX+k53gRPL2apRB/MayXAlBEXXvst1e3ALiXqbaWYRv7Sj5
128pTsN8X+/yS32BxDcPNa5k4xfP13p466dcFTglWy0xbr5ihfd68q1sZuH0N5+I
qRQitqFax+pJYrBaO4HCjYjeZ2nuptFMwnJIewoF6IFBjvXoNr0T6DD/z5iJGx1x
6KtTS9YOzv/ybznN76s2uYpaQKKVoVYBBoI22ZmAXB2BwL7dMh4JHVIke77JAFUQ
kw8SdUFF514F3DWLobUmkHvI6/OH5vTx3qFQaz+MEQpmAaHRyqvtHDgqnJc/tPNS
cydEHBZxabKntxv4HzEg1w8a7GgKRPUAacshyeVcS+y3TFuUB4WHoyxUvsumO7ab
fU45Sq5/hCD6jaxLQl52twZsl44HAIXJdycG/5ged7UNcLMTF+NlykVGD8huk9/O
A5GmScpLEM1W1YoxoKzQrs6e5wb51MkNsFus62GQ07khCt2xaoGBcp01MPWLOf6i
Ho3sGvBhjBAoN87+EeMTppjjs6yrdmVr8w7B6zp78ridF7PkKL8jIa/QJi6AZsLA
iDgdzEvQlquZwmZRNv1/MSPgizEeb3fSD4yU+qSKO+/ny5897vXGzlZlbA7KzHbv
B1scsBZZsbZLdx0wt/U3XBiahB7uOSzJz1I3iUea9bhZ2YTiITYpN16W4KxFawRt
atXHZTMtEAzwzDFx89kAcr3j+CBdrIWF5zTfQlBdOaaSvUhzaBzMxpBLMqkHwWJe
62FmT8HOphISa6vKz6Kxs+XDO/Qrxg5t6IHDFO4eKZKJMtSOM1vSmvzNvlkgfBWo
qlAx2Vep/dDZ4gLp7nY4I5hDB87Kz94ehkXDFNm3vz6EkymV4IUWz1sWFAn9vh6C
cl/KYtVvH+Wz3mroAHx1zLP/3Xx12Ilrqr+kXHNr7XtH2y65At4aJV+jyKDBbQZh
reB/UnixBxvvlxS7S3O7vKtA3u4UAzVlUn4pnDv9+TX+A5AeA3XwpnRDVGkMCTjT
CG4lYxFFx6rSHr5kbY9GBdcR4gL3gedBXDJyHrpanavtaIsp3kGDWV06waB7qulm
HtBA3tRaXW0SL9NmL18yDTlOlczQWMIvJfrag7IE7bj79QdFfaAzKwkWFVpy6+y1
/uDHT9EFXBNSgdPV05DabL/6H1juZlk60bm2aUsHECfBw1LsliZMtvlclLM8D47T
tPOyUF4VVzz00gA7sjF47cKNaAYCoKrNnsIcqjz1azWh6gCEkcNfgh/VzpM1TzIJ
GFqCY5n4KOxpYTlNoyWAchy0CW93ZsQgUQiexHbiYjisZCTgDJpTwzULPqYTUyOO
EToomCfM409OiWxU7PJkSEwkFt/khubo0wi/VjGlOLxTUWMG9Y09ziUhhByssQ+J
s1cXlFZ7P6emnkkU0XQE65T1NIhV8YAvlogsZ4cj610pxLjEV1kK5ttyJX9LRvN/
JGeKUMUMImZz11ATFzPT2eR1EUo/IZjajMbZuiLjr6EqPZF1WJpy8+9LK4+l1dKF
tOkAW6GLI0TbION/n15lfraTP0b34//zPcdN7QMuay5JFJ8qX9f3Mc8QupBNcBQr
r4fHuvLffFnzZSPlRK9aeNGdRqUVNoCWzrfoxwHOjF19tT/PAkqcV6EZAALvkVw7
Yj/V+OOebDE61mcJK/OBoym8mRaf0Jjgw1EecDxa6f5ApGKa8bm3jc7JC4yWZ8CP
Lxlyr336bVdo++Ql3/9u/xAVZukoB95oPEwUxuV4S7PyM3Wc1Fh6mqi0JH2N7Jes
f5Cf45nj5bwZY6sHpSgCezvhgGCxSF4heiYsd3cvnTGwASWQhlYn3fjkVVvqd+bD
WUHueII0esuhsQad0gHW5yafFybG96QzJMcOVIHTIR+TwykzK/hB5n3MyIOmK7/r
mNUw1rEWaAMoagi2Q5oem6yH52GJSqvG8MT6yQ0P4fprCGf7wokkVtVxzOd0TLvc
2MHYcYz806G37AwBZyuSQSeuGDmDYnVm/H7+1UXnDV8vqTeNLtB/hQmJAvFRU7FW
GJTMRja2UfOLRBCwfyut43wPuQib7K1Ky54PKjYmDrlbfhZxMxUDPzaPLUBs6s/Z
SMDMvidiBopszg7FQsfNDEz9GljLcDbakjUdbxeuA1Jk8X5m9O4VDZzE6FXRdQsZ
rB8MLeIAcsKSbBYHXb6bZ+DTraOWqHkpqxk42yag9tMOQG4EJyTrnbTsnTUyPenE
RTJVOd74hJnkXVFdZhUkvxQXHqMXzZ3tdoAucrf1CNUcJhGdBeHJa/QRNnI+h6Wk
aYsFH66w+9ZRZpnI82DSVBn6s8RoMK/wPGn7ctBJiLWsRCyeYjCOwhuqPRecrhRW
RR2jG5oi0tqRaS//Fnz49n3QpuzpwA0q2j4tERAeCkPSzKGsd19h7jvc8XU5LmKw
MSRbGyVOGp2Mf1UHcnWyxscYIEJOyRW1l5ixPGhikvI1Y6Jk6sLadGEqD/IAfBQ1
FvkSto8ajdBllEs9WhplL82VtFdYGZohFoRJ/G/ylr9oioNr9BkpfRK1UhzCLwIQ
DbeuCgaa2bFC5klI7ZBmBAaZtzMaQmhKAZ4vehi66RU3ARU+aE3ID8Ovj+JWeLYx
42Y+ZyPIpieU2xrQUqCbHUH633eILFYJItxtMwq7mmefm4xTclWHFBtZDqcA9g/z
lnZXE2kAEWQ3doKIqYmlYVZvCrngUxbV5IjsqwNpQqgloenkVmVA3uL6VBJbQEIM
Wi1XaLYyN6ZE/rYX9QrYqJAyer3sG+sQhMIAtUVFMa0J0alQtPx8bZIBthoRnqBj
ejkThkAtMLf3K1ErLQjE7kwgn7jeiI4ID1XRz47swgds6sR9p3gQfLGieyn++c4J
`pragma protect end_protected
