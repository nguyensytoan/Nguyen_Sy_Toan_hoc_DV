// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
um7gpadhPYWise4+WgWUYtSThwM8+hGIz4hE5cCsGplSgt4MmplbpjQ4Yxv8SmrRe5g2xy5Ty1eR
RNFuLkhBoa6XaceQgvsb1j0b+z8nO8+TUCJYttv0olvHPByXBYZGUjNpKz1KVXOc5KNyMv1kUbf2
wqTLD6ITvxQ2aS2EeSVTC3HWlIGI4gzBGIVK4+xye9RR8TbtwRbpzDAkwD6yj2NujB1ujQHWJwJS
zgxSCr3kzxre7TQn5UjPHWkpwpJevA9ZeCdgx3mDPdleixUaihBxm3L8exevXaxTp/qPGJHiUqaa
hLksuAYfOtoOc06sYJ19umc5Bxm6SKiebgcG2A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 30032)
tJrO/Tnb4EpsSqYs1tSGGjPgVBZMTH4ptcAcnw1/j7wa51T4MsG90H28jK7XzNfA80NgDqjJHidt
Jvoj5o7PM9s3YQ3ShfhG4sv4GWGlTrhLjwygEgCFJ4tqYMcf0V20eQfuWSs0KX/G3A5w+8dFwGY+
OltjqWAymgHcXXv89n6cFqe1ai3iwBSAj/O8RAX9ZNxU5iGp+MNYwNokilJbN37nCI9PQwaRChpK
VS+v9M/rN3e7MhBuGfAxO8cICFFnC8XLUwqcJFXyv5j9KZS0X6FGUcArO7tR6yuXdiGmtKAy6zms
pus7498jsrXHzqmpHX5Vhji9B+i23cqdti786vSXTnzMS139Ie5SVcT08gsSRFLZ58/wJQgVEir1
42NnJ9JidTpncjOx7Rs8q/PCxJlSkkSj6MiLRm9KrT95cdFOdHlftj3cjrSa+tiU+uD/K7h+N45K
masDfpcvm0BXWiLKn8c5jbv5kIm4eDBNm/z7BN4/ai3jz1GNyO29w5HyYeasQyw9tuCW9vzs8cR3
VuiXskRXnINBrAso0P4CudXiAXXWW3fQXaS3MC0nHyOPruYrC2jBUeE+wBMYVya6JmrtVjLIV6jM
VVYpi2jwWbBh4fyoF2HN3ArfFn9IYOzHjJMYHWoAAnGl8MmXWLmN/ML0T3Kc0LwaA6YCRvRd6uaQ
slgdG2nbSUfAK3svjCXQILbLMmUrZs6ucYcVRT77Bck6BOud0+aIX4tddirl8avvUtx1Ez1Ls7fl
IEl3xgbGVbbnAzJVsji1LpDZr6OQA4f/NKFOC5wwvK4/gZBKeJCYHBADQoka7AvHk0dtUAVLT23L
NjvCPD2Lt8goo88tX3MfyBv/Lh4Zsv23DcPApw9XbWbL9Clg+92MvVZdZj3NKjzxFjScFjtwFz+E
DPO06M/ww6SZU3yB0CI30lpfpEPhkSRi+f9rqxwzgrTUrKI2ccHLRR7e6eo2n+sc7sCQnfgJLYcy
tv3bbiurAb6NAWgmD1BYIil1YMkePfS6AlKzm4vN/6IKNYBHSfABHF8PrwNvr2ojzxDmAWl10Mo7
3BLfDltAJnSKm/T1GSSXuUEwBra7eyumFGxIhrjnk44U0gSfD95d7vJglQWnhcdDJGxXPPmToGh4
/ryUk5IYds8PY1IIbQJYv1tOHyxHKYPcz0VJEUsYQ6orF13GZyB8lj2ibh05xhikZnLD5ya6azCT
t6FBH6syxYX/5eqjUEGx3sI/7woz6sHegg64oI8U9j5iL5sQ9AMMdzTZwRGozj2K/pV65lHh7seB
IMuEb7mXUW8jDDYuYQkvgKb4hfthuuqs3zgYL/YxQNtmIIgY0mzNgC5bdkPnSmnv11dM13NfB7tf
xNlg86u/5ElC40czHdkfILkHFVv+g8poACy7H4y7p+eZc8yE3DmxhLQeQpOamW+zgMvGEatjoGAQ
4JLX0fBu6uCy4/mjBXs29966qnCvpitfeQxYZrnpi+mOcdPNK31mo+SBldXpZ8dRB4np6Mixl+a+
4jdWWSvR62db0xp2fqxhs2AyUSGfmeTv0FMyjWxPKPMeeQSkN57qNnxoHbw13qYgywPN/+TKiJi8
6G/McnheKcInkqZUttNq4u9WfY9wGS0Iv46hQgKCpkyQcG3UxghwEBsiyKdQNfvJ4qxzee4mobM2
zzB0aBJrxAbY4aGaSGHc7edTIR+JKSqR0eUtPCkExT/WPFUPLDfeVkUHZEs9gknYC6ZAfs/85qFI
cDpJoi0ohircLYNfxXZg6K595rBP9JJcJyPEQbvCBH5Grf8g1HYdPxiQfxJfBd2h+mclCqLz0MZK
IvPRhEEbafMvqDZUqvNaq78Boi+Ka47ty2S9Cjprqi6J0GrETGi4tOZcMqD7kqci59KS2sxGENWK
xtK4ORHL85K4BbCTBrXNmA58+OloLiyEbUjfiQ5OJmtHKxnHP7lIAmpS5snsF2H1XPLzX67Iezy0
xR4ZIn4g8OC2MhqN7uMOM4wwG8d+056x7r5Cm9dNgkh3x8cEd5xKrOStmQirgRtBa9mX+cM7J+eu
BOwlfxPTH0qu0Fc1uyFsPe93ooLsPD0WCOECZcW/64tOH1Q9Uj4nG6VTQExjmDtoyhATn6gxzprt
Xx79g4JqvK4j2zI5/yOmGPmw/Pa/LtpTldF9nej+myTXGNEdmsYdN1/UdztNt7jcDbfovaCUHFtj
m1qEPy0+zR/7qEa+DcRSHwDW9qH8HBlmjG4sRZflpLPDTd/9VBU9N88cn8FmZIDTbzmBZnCNkavs
fpOzEFb14qgibbYRWAcb4H42lXdwDlca145zj+BMNsi4mcUktnW/4lUvauNVRCFClCq5cbLrStdB
tCeMcbq+Z96eRspEYzAAel6+Rsthhl3c/h+BhIbapcqPAsMB7n/CHKHF1d35HOiTMvH5yscrkfad
XXtLuIqlvhqQr2m1PUSyw51GeAKe80YdsJrrmMMalt2KJjbT3DM2qW95ql/ZJJe0269td6F6zHYo
sH2/YUq8JP2v6i1txvhPQ1K7FxfJZvKqxMpeVQm0IThKC4q+BWNazK1hZ+n9L9V0n2fa1AdxDf5P
DqtWWpgKjMEmnkJHR4Ub3CIpLogTj8EKpFo6bFb2WncJLdLPaKANh/Mszu9vyBfYjb/odtOWkmYh
5bXEpHQsB5ix8o7lqgWLpTp+vPLz1K811BVfb8+OZCXvygmj3uE61EBGQVph5nXLxTWUlmadKGWi
JLMhyT9+kKXW+8y5L7Dtt8AjUOdnf0s3ZPYvWdXM5CBnHXyzpJSBdECFjRlDiT4BGWFTWXNrreW9
m/TNpEVDZFUCbLKbqNZFABJdZaJrQEzv00ITNdJ8OJonetRW+AupaMH2ogmJ1IckzHPM+H1vazaG
CC2SuOKDvTJ/WtR6xtsHZVALqrQE+NDevEsv5ysBq7VpmtiG4T37wYlW6yxOGH6fK+ja0qINYy7v
eI3Cq/MiS9c/P62zldPU4Nqy1V2ojvwcXb6+O3gNRZOU65m7Xv1IrZFqh9+QJKkSlETqKyUh0I7o
Zow6ebW2F12qKYj2EPfNIjHrLWq6etYayo0bBI10v4TUZHZM0jtRVOtsIFKep81Vt5Yfz7bv0FgQ
X9X0l/hUh8GLmttjXz+D8ogWkiFrxGcYBtXcrmdNM6eC/aQ8Ea5MNv7p3kNOtjoL3d/9FmdfsjB2
NMtdKnErXhqwjq9iiizU9UMhZ3/6v4PhlVZ3gXSjIG6/Op7EXCphyn2hGVsKQOGQuICAb/wCI4cF
etyEOExX4dIBkLYevCTo7L12kBd+6NbmQlwXv/4MGNlN/s+6LDOOZUvJiLeoT9NI6hP63axk4kxr
At89x2dA3I+3O5Nfxq4U0Ggzda/h00D+NBSvn7sGiRCITQ8Cka8/7JlYcwWBJbXNMbWnhNaXPzti
BzS/M8sAz7NY6Lx54IcEEt/dNdt6ThqmvwwTsJYMUgglHP4GNPvFHqWPxrfuoLETXAy+lw+RU65l
P3RkIQIF04+aXnoGYLmV6zkha5cPD2YwyX153d3gKnHYZBfQDkPMpK7/AD1vBmeobIlUQ/TtBKnL
6KOtZ+4i4L/dueaI2Qn/JYd3EZWczFoyz5sR8q4HSFS6cfjPo/EtVHH803gRpTdEg2q6iOPY1LZl
egkYwh+qqeOwyFV50uGqMKFZdDISMcrpJ2Knk90dMUOrWbnNEZ0217pWcHIxDPeA3g4afExB+sB1
gwzbE+x2P8TF76aMgk/Eqs5jM1yJr1av/N7jSn/ARYQn3i6VbmI1Jj6WyxzZnzKh0g8LOxu/kTnU
eEIqYtprbymfZIAG1lFH5e0neqo0CyylhZE5geb3PTh+UkugAXQ7kwTs26X3s4CRoB91v1GcTKj1
IjLoOdz491vAwIDMqxmYKMb6xPNILHWwhXYNIhn6HfQ0jmPuMnlZsPNPETcfDxMuzKJd52uQBKb3
ykCV2Xy7b92jgjqD8Y8DYz1giB8ToaN1yTR9ykSgctV6djlaEctwDjLXdDwCRFL0BGGnom9flhje
CRXowZacGK+d3/MzZ5CxT4lTsF1lUG6Jh8JULMQoDBGjFpNuPWOfQMBvXL/MUWBlQlGz+GTD4yO5
iWmqwget6llvqAptHbkTD0XW9RuqByVifBNrwrDP8NgSZ8Yyn6yflJOKJvP3ei01eSlV338NikrF
uoXTNuyesGSgiTYncLbtadhxWiYsiELxbHe4Pr5E7bFF/DGVcRJNqZ/tSBSR2ZEmBeAZ1Te+3Zr2
tqNPZ5bgwHE1mn61qAnj3dJ8qhpHHJ9/RipX9rF6RLCPw3c5KfM9RG4SVE2r2pCXze5jjHmHXTFk
dnGb3qOuUXUIxjdM/4fDSQXgFJ7Ah8cZjznL7a7DBxNJ6z6jIRZRIUKrFnTb848sFTDUpwpCKrNW
hOGdSXXebBZcud+hvTM4HWSr5V6ihLcS0T0j9p21KxpM0pl076fsSqbD+mI1S5PmPWGsfcZIrNTu
OxwtbqFWxjZrPQktTWnlr5aAW0uMymk+xe5bByJBNeAgLnevctqPuuXwflWm0L8mgbVfjJO4u3AK
J2tqU1e73802h6n3GYE4zyHz1c/qXjpWQ6bhZWmEH2EsEl9LRk/dodi1wCFM3moOZ2lBFLnEfhJy
bpgY0OwvPdj/GtIMwN4HYhb37PX9RYKiDbq8Pwor1KIq2XtKrqTyHfKBBS36KlRADWUayFOXmLF8
r+Li7MzNfEo8Io+LS5DE0ul+/kO/fFE+5ozNZ3SGt5luuAsxrbqje4IQz6Wi0NuhBUpcLT4ZnVb8
BDSDa33ZiqCMNLVkt7FAvLs/rN2GTEFhf69iVaue/KqztjwIpXhcbxbCBZbUv3xXhqY0W4gEpD2W
RZFlx1VOjQcFd7JR5LM23H53taEaCr7A+TNuox7/MxGtlZFPwNk2/O8Pe9KKon5Jzcs9M94d8ZPM
IJbosXWoE/IcuoLByp2xRjPJdtmxOlzY5dzdyXlJS7Mh7GSdxy62QyI12l0KV6Q8LZzW7tCsKcx+
I5YLolM4lmhOM6o5rsTIMr7ZxUt79TxxeMC6L30H3ioQxhfjTVmwXjUZJu1LCqRGucw5apPEJqzd
YEEz96cpMGuDS/mEwgXM1q3YxB3+Pa7v7w7tdzKNkK6XGs/1GIATL70Xv48bbLQCYO2y0Z9/xu1I
iGZXPzoFGGLe7gwAC1ZnTiEUNCGbDQNidsKhhbMnPcA4W3ecIUj+Ue0dTcHLb6GSdxJLWqI0Uygp
jIAZQ4zawvKNCECw+W1TyT187pqp+ZSzcWm02NplgfVLgvaWIHHXHx25xajmPBcKJyxJFYUUd/11
Takyc+jJCMzvRmqhoWqTsf700IAbxFWmO0Ei2SliX3KuSKkavsH/p5F09FMdvftU4CU8+mQSKEuk
rZcAxp3O0zKY/wNSXmw5Rd7DJYK9gLkNDQT6EGZ1fwAIZTCM3tdjvwlgEPXFK25568xasdDwa5ZI
jAv5kIqQZwx3ZSgnvO9piDd6+ECYqZw0xqJNkjlPTLebyl9+8lY8oWeFHhDTrYh3YpJ9acjfxUew
4euVyQoRoGi8SgAfn+Tt/Ddg1dcYnQEIHS34dQbFnHumECxVCnQ2TPWvIv6svBuIm6dcb8q8EyqQ
VRxNkkqqXM3UrILjy8J/T/Bx90WinBBPNS6PrMKM8LPp63pcGw8kO4PLMWo/NpAHbYq295wa7p68
v502KTUKx81yBJK17jb4HEERwEn8LYqiWxwl++Lh3c2bb6LgufWLWXFzxJgbsKGy7Z2uYsqeEZoH
UstV1mjHmxyqWxKnqe/kBXPraRVM/bhigaF8AKmiOwM+5L8eiFtjKoNYVR7p3bgV/Ivqqp7bLDLJ
OD6tCJZdp+QpDLqpyACt/4Sio6xrK1P3XQKa7fHIo0YDHIECMx4FdKy2g9/BFpV9/NY1XD8UZvuo
0aFDKHty3MVFr11Gety7LVUsaS8fJ0okeqqZ2gfSU7S/JR1uyIKB98wBwyNY2aouO2dXNi+9DrmT
hC8Ox9x8I/1MEHn2UQxhWg+g6MVkZ6SF9pAEbb252V0PBVdoqKz55StrFvLyizyL5QXtlYhQtVg0
z5csVXgPj+mCZNhUa6kk0zqFP+k8Oy5m4Po9RJcWVvy4wMsg6jrd/AS+eOQSNUh3tdlXcfmVbZOq
uyUvBzO6uG20MKBH6noUCIeZatlc96ng+WnoKP+koCS8SSSXty8VWHQ24ZY9smb3vInkv2ouAkfb
yuvjz2EpDQbUTmUWJu0a6TIssrejA1JEntucA0OX0vjCoy59aZuOZ/eU7Q5Oib5XuHAUjjuJDgeS
26yr6Y2RjYL56dHgU+09FPQycDQ3WjyADpJHxISjuuGr6d/xl4a1maH7hTbOk0RAVrDB7mD4kgwE
axTyUiLN0KG2Pu5+euhCPfKkcQLWr+dyBxOvl1PaBSh2uhY73piBjzF+g4coce37vbKI8Bp1gtKF
k54euwNMhvqDm31HrFWloX5ARlEHbfV+57tRkJPLpEhZ5Hh4eJOwCzz/1KcKn+jSbtm2mqGOrVV4
ElwZvFYH0B0hAyzCyitkNLtlfunv++x/Pha2rb8HAv0Mxc4OXKeT+Y2kREHbNHBp+2AQhWM/PIWF
cWf20q2Jg8o4aYqDVymbKjdxlIbVvf4OfBhc3BFvm9a726E0bZ5bkvbZD8H3kqzoZ6VBJxBZU1CI
EdoLisQhTTbLEBbMBVRmjbp8K/HHvoTD6twWD6TMeMtrGx0ir1KqH/wvIkU8wh47KWSzeHnm20GZ
9YyRKvRzRrHYeyZqVuXaDt09vCK3XNjxVm/zclCJokHDPJD41gx7FPkeBpNZW1xPCW+MlPbdNdqU
BrTCShYjq2jI7/YapLPYxoMnBffASa6o6FVH4HepO9CtPRFzYjbsRQSaPxOOjdxEzzVNnmb8HiEx
1XPMEA2g1Uzfc6hHaSEjrP+/D2EURPgonxXzZcceIpXzO0IfXE/PNmHHYdUpkgl1yKuUVBUTCSWW
WxWu2gfMPg2buRVcQnuyhztvMlwwVpoEW6ZhFY98Qrv2rPjAqxx9cTy4UfjYitjvOJHSL9Ei1og+
ToOVofC5hALvCIrXD+uoI8m5Yq9gNb0wT/N5NbedhqpMnkkGss8/h/baaFDzJL25Wbowrw1VIBWM
OSgs2V8uAv3doJjSBI7wFu30kl7Fy5n1iMY0BSgDlap/MWzq7gyQjmYduQjwbmVMfrIYdZ+1zmW/
6OiAUO+KQ8U4t0l7v8Qde/LI03EnOozPJvQPcrV6INPK9vxZgVOX1vhvGiFAVgNUy/NI+8D9QGZt
WOi1ei6pZcq7BCTYuOtIfgPRdvw+ZZ7j72gOsK6fJns19TgRdpbZ4/LErM/2+SQLBz5btXURlA5o
ObZXQxEyU8tUfOFI2oLsXchGNE2Lr0x1PH8QXT36O5V1x75d7SyAE6dT3qV/W1EeGyGSLEALauKX
uPCe6K5MvRVK+hI6VtzU3eRXp+L+AYdlHNipq65MvebJGPO1O0/fbPNfRtIK+YbXqOT2rPgR4d+3
NKKci3iRb2kCfvetSE5U0ggs20QpQh38XCdb/iWz6yeOOHdEzWN6xOJBP7A5++Ojct/Pj/s+/5SV
QBt1zHyVzjTaSXrS5z9d/VdF89pT38804lOeVvlWNviVAUklg8KIysolcznzSZXXugpoqVmSHagf
TQL5bz8YOxfkjib9Lk8Pg9M693+jvyDg84orvecXsWqAgFhIpgyaN7SACt8J2X4HphfbmUrvyks3
s7/JR6CWLlo6Z9qcv0vZurGes39Zb2HM/B6fbuvu3zKo0TxrTL6nwHPYauagrDTaekAHQUb1wzAq
0g+n3pmEeO/+eNLb/h3O7QSZQxVMjZp3nzWki/J9JCOmgoCiw3ZvQY3V6/jEBei9eyYOz6zTTJui
EJRPxfLB+uyf6hkUB/enkcsnPvFpnXO4OIsDpKYVDi5h5fT5vLRprgavE/II0GhrhOTDQkVG0Aqo
/Y/d8FDkcQN/dexoPKa1WlzGltbL+gtABnSFVcsLynBD8wCjA6f+MhZ8ec7wEKo4uNjLql50flPM
D/ozaX1PMsGczw46dnTvly8KDDOyaYg47/BrUihbysWGtVrERQqtx3s0+yqKCw8Aip1PReXcIOb/
xTxT1WaW58YMoBBWFRCynjgLTxBv77L5T4z8UlFt0pqYCTQ4z1TYxTZqr6EpwA62bvRmQIz6nP3F
vcnMXXo+kVUmBgNZ21XTjXyCbaY6Vh6Yqkxro06Nh1QteAAx1IPJcfmVQPVc6UMpwGGEc3kA5fbH
Sf2nsQPuX3kqDlIE/V3tLb0pyWk36MSSaQVePgWI8njp2/nM97ZlZ20MVh3PneJmFyZ3unpA9eUZ
5fEoNMsKP71i7TysCxaIFOKt5UiZ5LZQMd9hwe4Mtuee/8qxca5PukBJvUC5Tu5QCoPujYuSEhqi
XPk5ZWOPx/EUPYp4chCbZPJkdDmsE67diUTtOvvnUXUOhvsM6ezw00FmUwDnN3Dne3thG7ebHnH3
cB4beBBxqiNXWI1MgiIWNkVhg0wQVxwZz1AU9zTEWXtSV4JmYJgh/QxgkKrMX1XLBX4JAE2yX0EF
CPyp1qAJAOxPu14zwqjQksrP+6UPsXpfNhH+xKDdW8SjWPtBBDjTB/WJpEMx9eVpfCiSYqWIxftt
kTXAFRFDOGL0vq1zekmD3lazW6ArO3p12igCR0OA6f12HRAMJLWyBHx/oPGR9mqSa+8SRC8hb23I
+dSPOh0oLQlFnbrjJt3mFOmhK5MorCD2XoVgtbK2LOxmz9uY8oqBecSjp1Mekwo7K6cv3gqbazxn
VpZ1Aq1Ujs2Avtz9UYORu9MzdbKPnBb/9nD12FXNjLKG7uFG04DRhgaZGjqnf+jtIPsLHdtUhbr2
ibH314aXJK1c4guU74HOBrSJE72JYU+Hi+Z4SLcW9zD+QxGolb1jZvAahgk7TUWjC4lnQ5K5J7GW
TuWtUVQDJ+uoPuqPVrkFC3yUgKzanOR6GSDdvj466oWxGf66vDm9uKNlzp+3RqV08ciiiYUw5Ijf
Oz70dPlfGHHIfwu9qrpkc2hr1u4F38bpEr55Gfh4W9zOwstamU8L8uzDYx5dlzT4mFGR69rC50QL
vQc9ibIzvq0NnVtCrtyTrrfjoPQWCMmUP5cJ19Js6MT/mNfyFIgZt7EdpQcW7V3NfcGH7K5i+Sfc
w9oOnWfk+zcKZZH22vj39Cwmoucdc1/87K7DEVcVvqDm84S8VNidKuselZ3/dEPQXP15gOdbnyYx
rurlWFUOGF8GD3s7bIl4gEqMbOeMTRWFDxZEBVETjEVdzDYjteBomLXG1t65o/oLx4c3Ew7wVrgp
Ddb7AR66tkI3Sy+o0Gk8CFl73xwhYzJGgeKH1g1IID/oh+6mSbnTmYN/pMD4iz7LUp0zkso6ORzl
mC70u2y9a32zIQFqbMIVzjh78OKOUHpxa+2oCLjrWyQ/3573kXPfZvtz2AwlYSCZBVWyaVBSMff6
QsaUimdwnSWKgTHpAn8ba6XRG7j5VxlQSFkHMNsrHCIoqyXrhJbF3TP1oq9CCeQcxcrgglEyhjZ2
LGq7SljpEBVsCpgZiW+nncA3BYN+1E14SsOL4L034c6KRIffNLmjOQsqEN1JSMXP6yVlI9w3CiHt
Rx0lkOUhfKbPmobKJiAoDu04inCkRgFcVjhgzl9qKxOrjAkPbfS57C4rh4fP7Kl/Bc9whYpm7rLp
Wp35e/A2cnQ1UlvG/MD/YFOBjBoKUXOMV2fK43DuBK3Ff0Gk5Bt6I4kvTCv8E7wux+LDommG0PsM
0jaYOOCNloqGcYUDmbMLUQRzfngs/MipEUYwLU14RBfphS1ej1eNkdKWoeKJmyFect31npQPCrAC
o7xuF5Slnb0yMW9RtA4vr5kTp8SsVJKvvXhRXyi0movbxvoU2+yKdSFPeb3JgzYSOBGEm+VfyDIL
C/MT4rJYccMfauvplBbuYGzpZ2fPMeaPx2ZVulUEHu4XsSTxn+8ZvHdKyjzCoYcjdw1IJG5+sHqM
BRY1YYmIvY7KPkM4GfwEvUfSmQb/yUzilY1OLoS7GYB7/9uPfmNGgF/RWdpWnOwMRonu5PeB3+B6
SJVDGvHCJJvURrPI+SGDf8xw3enOxw3iy4BEwPCqvjaQW3/MgTJ/GKZPB3TwhWdfaf4+03tqL2S7
UrXFPdAlFPKf47e2FldyM1IqRTCRc1ImQruRFwF0qjtIUBCgGP/hY4J894+Ci02c1fRGvdWt5FdG
32wa6hccVXLDdOnfBw74VWx+dU7IFaVN4IbJbNEUFp2UdwFH/eZ4km3A5hj3kiXwW/kOTIa9YeAV
6FZZuRjn5jgtNWAu2GLwbBFOv5QuEQx/K+JNyRzU7aGx7Kr4SrKCc9Ha1060MFyq1GSKh4Ka6AuB
Qy2h47LDNGPKS0xtY1KUVDOe0ox+usks074egwwAtlvYiq5zN0PaqOkZ5R7ygfMU1oNvrdt0yq4G
SVGFB99oOBB++wbXvxw6Jgy1SO+oksNPgWEgNr8jALUz4OKFNGdW1lsepr7dKLGUAS43bw3e3qes
ixb1rViafFChMHyW9gmwFxwkzTmf+Y24ITjX8lNTlBAmwvjhlTpBjka5U5VZh72C2uT/86mjznw8
Bohk/kNRw52o8lknP00KvzG9xuOQuf9tj44pno/BTRiGxNqwqWZZqmExOHz8EC60kDIP6wb3LbEO
qJ978H2VNLdXLVjmIk2ADLxovIPKRRFHG2m8rCQ4LD8va95vBpgdVjw8iszPPAewOCma3egfcGXv
KS//Od1TWUb9w/n0fXJ1B7oBcRaMllw0Ds0yEo1zrgnoTPbZeuL5vXMNFWAlQEmA/PpEGvlLdQM7
pwSla3SVmwVFBxuSvcHh7486GccK7c1GRJ31Tfl+cvrvYScJQyORreERNcT53Me2iZphvPxgqUcm
mXSTmiORcTCu++wv+Hbo3SVmEey0z4B23Vtf3BFsX9nVhjOC2wcclhGpR9jTSzCwuDHM+N3HUK96
kLWDfA2nG8UUtUtdGGFL1pRI82fvPXZzlykp0iH4MCWHKQSWPm2fMTZ57PKkjV2efrcT8ENJOXdy
s+F4quzrfvfhM5On8tmG7OWJYEtU5O9q2IE0UqswH9TbPj2IICKKAHtf5u7OqN0vYSU+gcyfySRm
3DyBc/X10iLvgyABVqpSkabQXiVo9LEpAekUqcoouetgvOxUMb+aEXrAcpm4Z63M2SkO6YxvHxWr
X/EbRzV9MEbqnfyJu/3mJ5wDUpmJtgMWoP9CUWlZDNcxpXf/4FF1yg4QO2q6WJs7BiuMteRgmtiT
nXtyLepNeCGGpE7M5lH+tMWDFG58krrcchn+kwLgNBPWbzZ5g+4TcB54m5a0udkSH61VI6Disd+U
r/7zGdzpMezQcIq3SSXoF96XbooMbhsZKUw19t/3DKF4Y812YnPSMw01r/wi+PFGFr+tulVg1P0I
0FrLma7i4dg8FhWWcR/HKsi+Bv4mSK8mpc1xZVrlKy3LxJMFeY0gFj0J+5zVVI/AQB79vcssQRcq
O837Ec6PIjgV23qnE4aXwQHcjwnm+WBDo9kHAigjnsc4vQt6prsYf9NfN3H7MJlKYug7nJhxK13o
d8HMyfKlNjEGNYkDaZFPKKWsrNXQEz0nOxOObLc8y7yvgQsWyIi09yYZJwrFg7wwWlBo1Fn13sj+
DF/4iWyQ8NnUAxmoeuUzw4T+nwbpmp+TNgGIn7O0CHObRkzTgZxeZpF9PB5NqTvIXcfI/q7R7WJN
maKiNWpJ9tnE1e3H37f2Lw3WAR3Nb47l1NRJ0yEzB1jirAYKweLJ832yr2fIJuO8AeCe/MP0CCnI
32/a7i5boIHHYa8I3tf0ZWCdJavQF8o2v6e0oBJpe/rrr/Ymn7tluA3Lmwujk40KPk+Dgcqk8v4p
vqZW7d3ThVH6sM4cxfnBkaaMNA3sPs534jBHcYO32luGzTcaSdVvmaGIco+/5tcb7iWbI1bR1OLG
uKWwMSQlhEukHmteysyQlBL6mz0lHQIv94+m/20WhYvPYwQYOzv+09YJq3BvgLdbcpo8iljid30x
EDbpTY60VRw3v4P9DiTvD59/+Uss5eW+TWcX5UAg61CsnVAWqMMIFokm+2sGU/v3O5e7HUBc/3N7
nmK5S9kG5wkYGSl155hpXrro1bOcHYaRSDLaDuSh+CEOAMFagIX+/JWkvxrt954CT6Rn5REaw8t1
7JY/LOf6LwB6SZwRFgs5XMH4Bmv1NewZntufVyYyip/dg+tupBLN3VBpcpwMXHP4GZfHdFjL3CQh
n4rGtXFuG/iZ2B3Tv0T5JSZRtJ1B61Fb27DsGECufnGDl2W2xu+WolbDjAj4ETxZQ8X/BzLcY6Wf
tR1pzzdNGNBQNScWdpwET/RTnYurU3ptIXnKLY8obFavu/4KBPyW7wFeUaTb7+lRaFJe9srW2i+a
KK3sdDg9GXrd86GwTBqx2yJCC1bB/ROTUd+1n58hIZ90tWlu5BV38R2FABvBt7FQRtqQ1Cr2dxkp
yHPZALudYINohHeUBEnh7/bzis6hTFoqVgqCTt8FPmS7lC5HDdotYZ6P6Ql8wkgN5aDo6mBh0b9i
UWfqlbNihfJLJ46+gBQomqs+WY4jldo7dGtMcH1i0U9rafglQwQv6q0YoXcjDPMVmsGNAtlsHyLc
m9vt6Ri5gtGcNNaQpObXKwE9XCabF8tTZasGAxfeOKPxV1yzylqDMdrbKmhdaEbgQ/US3Ebh8Yey
Kmh671EmHokgDeKD62S827xAPk5BhbJpLQKtPj8Yb7Tf3vIoI5al9XSoWix1ATaEgZkXenYpY1hw
H04S1fYVL8RlAklB1+Lq6KtaVM/snAV76N/IwN3OxS5Dhrn6Y9P2BHHLYsIDZI77z0uEJKF6Kq++
ldgsFfk9yZ7feQisjtHy/phqXNMqu02auHwrlwUzrj36z8niStvzEhDB+aoCb5nw3X5SdGvWMJxf
pST4kZ+Dc77018+9W0vQfgxZ6cNhFQd5uBJyIW8/vDDoKp8ON9t+59z9laOZEirtQWQ3wAdzcUwX
W6/HJGrV9tx+/ZFfGXxhZuaFwJ24WPJzY0MqwhXzKutY3AxaOQ5Pnsq2Qr50Epr+1t7MHZ31r/8m
l8qa07xvAAGol2sxFy63fJQpV51qKMRMdedM29yne/T5Fz98+E8Pv1iozhzmtSWYmGo48JJ0b6FY
rNxUSOtmkhuwnKH6mQzxaW6DvR0/nxXWDkbm1FeZkqeOOLvGOiF9KBFdIHNZ3hZinvowHx3RS8xx
3E+/EPDfc6dxM8K9RHqqshZbe6kFVBaGpdslq9QiB3V6h2jEu01zsA7is9WRVrHcgMoCeXi1PE2/
qh7iK1zTNPTomjmETwEq3Kg8ifsfyJx+Ztf9UP6Lbc75tfk0S/VjwH0efugOP66mp+np6dK7fQu/
UZJ6gLrShVxNCNk5WJ3OJvKJEn3OqvdWK6mBsr/1JBeSg77Dex2YvV21Zzvj+49u6KRcXE68Qd9D
+zzeiN78+cgMoXeluGwODiqF3K3NJfxKxSXrs5Zqt3Vrr4wr1hkV3CCo4XLLD441FA7YqtbUvTsp
pLn8aaFguMrJe+3J0SqzeFzqzvtg/iDP3blsEuBWXARduV5VnRb9Pj7IHpjI+jimNPKnR+siM5Es
crheuiackjVkkP3p/82wd4sqqHsgruKPPImydBrkGnSQVv/FQkXkJmwLclv6p/QWcWevAlIzfOA7
kXCryDyF1StEyqWyNjqbAvk8qa4ezzC7M81VR8POJaREqc2rLFZSrhgwKVdtNe5vX0VKfB9+qMc4
VgW/dNc2Oe/7TJHMzZGTC/kGso6JDa4GZH/t8QqUboRCc2YuHZOy8OL2UX0T1lH6H1kxvXzP/dvd
vCbPE1wdifPSI/wUzMAsiVYcoEN717qokHM17BDh2B5pT9O99uJBLH/pKy264gPR/nXdO0TYiiOQ
WkVL3CU/AwOHYODw23xYYO2Ikfc5XhWpis8BaRlg5QRQ55AyrLvoJ1OyBeKG9ynwXqa9TuZunp9B
WXz6GEZqWsdUORsp7gJrbAxP+E9VeZGu669n/E6m4sY3djK4BsYCntAW/wx+lgssmkgSQ62jm3x0
pq7xYhePLECLB53X+E6mFJDoKkJ19zo0iLEh6o7Lse8pN1dbRFJ8s+7sPO2ZedOTKYQ7EWurEGkL
gd5JXDNXehSm/oLDZTk3limeuypeD9wdMLrxLaPoHUEJ9KkxOZbp3LXzO73CKuO4DRf5mQ/dqMJR
IZdouWX+vJTBFTFMb4xky1OGrjwkTllH+pE+RhkgrgzzgkE+R2wJ1kqNRbuKCKaHuP+Yq1yoTFpa
VpFo2xrBGs3hw/pWF/jvn1kJu7gbHz/Y9Ec7I2kLW153IpJaEOBccAFewpamrgoYLw+Kzo1mSWcR
hsC1AUMBNLSQ8mVShlMgzz1UvTq811dmBUmBWPyWlfljtm3D2eHYHUmKyMXJps1j00xQFBggeXFJ
XsoxlHCC8oDREfqC1am2MdNLyVCMeqc6oelhDCkOalRdgdSr3omintFofl0JozepVBzPBbucXb4W
v7jA0Aq2C3aCXK4WyDRF/rSwVRGKkX4Ubg7guWDzrcymfwgUES5HvsUJkArubEty/sGVb5h9Hhim
BHXtYT+ShPYWbIIl9zTSEMjupJBcpuJoFuCUM9HJFLmnnQKvFVgHuoLGlYE/ov5H3nW4y+XBqR8l
Lc72ioqUiWL7lkx9f2U8K86OMj52C/5nMCQx6OG0mED1tbyODLgT5JU8FBL8XrWEzgo09H4nLfHm
U4Joq3hpL+MOq5JccfwCwTRLXmnqfyAxlS8ETE6+SNoq5uM98070Efcbv4GP4LmGsRTiLKwQP7wt
QhcerIU/RA/CIT6TX6m6TNF9UXfi9pKBJsEVuHLk9tz0KP4nb0F/gonzqhUakAr6Dx28SyYl1PS5
b0uJP+cyhnXkxnts0UVS8FRgy/Ku7HmNHlG0SH7kIb+kWv4BMkiW/eASSxCdktX7UVtOk+8Dhwls
SmdSLePW32CXw+BGSuoI1tq7WlJX9xoJGNsQB1iFkV8vwUACZ7cZuBHQG/B2tMJ40FEeq9+ZTkkL
KLU1F7YGtEoSKFNAvO6KWdoMx3ZwacpdlmFC82obCTqOsSvyHwbHMOZRuEBvgZtLrJmpG0+JBAJ7
cacoc6Gf9yMPAnKZtRvyIvb/fXoLxO+TXOCvzjz+LA7HPQ0NNMZObN27BcJp4x2J9A7b67pVT+UL
yMjcZNyBr1lDOBmjHu2IZn+9jetpwlor0YLt8hP43OQebMhh9SacM/ZC59QeC40OWSYRz9ZUmhR+
vA7yUjlzw9cQql6uz3ylcrPd1hs7sHwxyWYYpEyK5lgsE5197lopWnNnJLlfLNtBMZgCKp6B0PiF
csmhSxWcsxZKra0F7LW1TK64lvOk6QIYtCX6BcI/ByjEGLvg6RBUGY1Av3s3W0/uSAYQSjwdeB1h
/NZmc2RqVLh6pLixaPhAL6tkQ4VmZ9acosICt+b0174cPANNvMmotRl1qKT83BZa7XqfSl0C62JK
Kg5wEAU5H6+H90IpcQJnyxJ8v2Rl0zPZAOrieAtZt1UfykylmjgzbumTctgVMkTkKnT4VrTt0Ts2
wPcJwe5sfDpBIF94gYPDs2Q0/2Fj0xh0bXbwRuRQdY8qI2j/ffNSI+hihbNV3fe6z1xawfMa52yj
yTkeUrBgJgpMefwGxjPQhgaf52MIpLfzD/lb8gXVWoigA4GvgYBNfZn05XPYDsFm7DsIxLQ0DpTK
H6qlmjvIhzHVfB+SLssGo59+q5fX8w0Sb1MQiVFb60bs7gFcIaDA/jShVtMrlvN4GDgbd1dw5oiR
YAhyrvv8wPjVYLUk9tfbSjFIZyyT8pNhp87dIuBFsVRkP3n7Ee2g6oxYuNESX3bBTNgav2E8zTvd
uQFgT1ek5CMUXa52G3wuSeUeT7xr9NLQRnIJEjRGu3kSyaPjwXz4tsnMngByuc04jTzsIcmUxr03
tTymG5SlPX0efzLfwS40Hp1zZT5kIIAZyf06Q78bwwTxWHuMZpBWwoaBTXKWymkqN011US7tA0Tw
VY8Ldwyyir6+Vqldnt8p96pf3oYh+RHC0YM6iugQwR/Dmip6XUfMwYk7nfK4CGEE8aFWCyRceJJb
71siNeSkj/VQGuWIQjbh8gDAZ+QwOGJgstz867LvOcgcziBzsM/VW4cNAHyQSWYEs+RBHCJRspU1
uRwRXP7GKItgA3aaDrGfQ/z7utdEiVyg3kEO/cy9555rfdd0R0vtGrt2pKK0luNyj2Fa+wj8Vqq2
kvl14zOAChqCerIpCyQJXW8bs/FTltIqIjpbU+z3h8VkxlqVKxFQsvEunX9coM3r9A/i+GgNoz/T
rZHXV3JgX3nnzJ6n/hIwNn0Zkh0pcHs76iI6CY1UdGTLpOq9K9C1VlkHGn7+qHTF7rovr98MLgSM
0jvIiPUf3XvlechRFFXFi8t0zcU4rsD+lCrviM1zqR0ffg5/ZjPHjKBKVr2UNeA+ZDjxeTSCo8YA
2ogFHO+4590MZW0FTcsrA0T9mSI8qgr0PvjjXaInWN0sBueb/s5PC7HMH5eIKJ/U0ohz4Hw0/IGa
lLnxdcykkWoO/HJFnqQwF7WKgGR1L83XvbTmMtTsw/X2Geo3KnwAWpDfDueRb6PPjuTtB2LgRyPc
uCfW5YFyW6GnacurV58qKjxX2TNRfAchxm5b/mu7/UcjKPzyCy115yzXZBc+mwHgPt+oqBNM4OSY
kSmDMjO/ONyv2EyYqkMAFvi5smcgbnq5zE1jc8vy0AqJmyplF7Lp/4wST77Xvw630kpmPpWFDRKm
bW4sWlN7T+6TCTkYyrRazphIn7kBI6eXaW+mobWj8wb+fz+c9fIUY1nz7hjm5cXReFQYu2EkNoMc
NR1vvt+yjzH7iZy+icweWUTqXaEvrmdScAsk3zd7NcmR5IHodEe32gj8idTNUE1cw0WruqwiEPGt
J1ce8SDScf668LOLyMKi3pwTduA5uxXzyy6SsJnhO6zVk5lwrtvU5w9qtzsvLJwIfQ5rBNpU4Ehu
MyaReJJHhwxZqQt2lCV0VCHo11uJ7eeCttxneJfjTwn4EKkFCGaLvMPrcR/mRBD4JUKHWART7f4l
9QG0zvB/RR6LdB9ccbbKAIk+W/MCEX7ivGW3Wov3l3UV4o6PDzemeMpAudAFowq0OJn2WUBm4XCd
ocsdHRl8O0b/vCD8Vx4dsIXdLuAyQEhyFz0xzrpX3JOqVCaOTsgasLcNE/za94WroIOCxyq3oteX
3ZPEwcRwjcX91btzNnNukUr4gcOzlgg0Au68EYsT5DPUAgjDHnbG5jLBca7cWk0coNtYPxD0KRDM
1h7x/7sJ/iVK0SMSMzg9uV6LBaHCmhyaJyX0m5m51krbytrsdwS9fgd33X1pYALvW0EIm/6wafKi
PdwmRbS4NQlPoKxRLcXbUVdYyTHl6XoPS1gfaFx33ov2zmpKz/TSPU9z4FrFWnxSMYtHNuPML3aO
JXR6/jTZeIMqsFki3Tv1Jg0FahK2CoMMj06vqHPy1dNjriBpu9cDHSUXfyMAkT/l4jkP7gD3Ulub
fEH/MjzCOEK88ZuS2D8Aq2rr4Co+dKs7EndL2Rz77b0hS4U+3gmNq01duQZrRP3oRAkSiKUs8omW
1G129zM97zkCY7EgibPIqkN3KnLDheq0GvBnI/EAPMvEZBnKdW0W2dieYzf5MYRXfr3DLBgzsxJX
QUaTBN9IGhH9Mh4qw1tdT/S9zg75RnlDr9T6phCyJSvftKehUKRQ8i+Yo6G78j3sDSW7CYNb8yvz
d5CIMoGE9vtLzPs8O8NK8eKu5MpfY0Jvh1ULsDUZMa48/4OXD807izPBCl97+1HcaFf2AE156MFZ
/6ah4csqGkA2cw1eCmTg03L2nYWrX3mqMdu5CEOseuZI9w3DfJYp+sqmBcoWUaEBxkK2KQSxReF9
dDtM/mpRW7KWSlPYEEEAFsrmDK5wH+sP+iocPQPt2r8KM7BLRAfHZeov6ox2CEaGDYSXQLwKKNp5
3q9bnodD0I8dJtJBFIJ5K0SCGWcoys3pGnPMhsbwYzxqgRWo092kTi5o3sT7wYTwU4tCnOomhpSB
que7zxToN6CAarx2Bu62u5MSuhO4O9bdljOB0anHbUw/vtpACFCDYnB5zkvBQOiOr1uPosImd5eU
wwelbiHcECYxqjlUR7wVJJdwD0qJBTl60xhXmLSQn3qxH2tYQkAaGQevj031yHimIIx2bgBe5bVu
ZNO7RJ6o+rQE71uh+uZ2GgUr58ABIko7vNnJYWpRnywHbTSDRZJPIReqhYDHijTbd9VzuVTykGtG
R/dkHXtdtZhv77WluNCV5u5bHHDD0INxDgv6byIkGAamN6o/uZ0BFaMarttFUzPw+QjfOETaX4Tp
gEqmRWZEv0ICZO3p4uAOEJxBkBQ0sT4C5eS27IA6S0pSGmEQVVseolJc3Eoi9bwRZ5jAD/Tu4bHj
96+nzE1eJoqLbs+FHrWfHPreFF3G0FNEmjW4eL+6LsjG/QN5kXauRICZTdWXRd18Q0ZBTJQECZFR
SCtIgLaVdpaiHfwNVlM1Zi+2bvskCdeH6dyr8VHxqMmUr38/+ta+UcXMzbyMSDPesYYQW6j78wzk
wvB5IRvvExRUOZTey8CgQN7vPmu30W8uJsSczXWKvHa7gpps28+MBYE99yQTffT+vCu2fJZ6YTOx
LxBoBhZf3Yo6bnLmvjsPVRBTVVLVIQALj0QB8YNi3tfnxuN9B5SfJJPFeJ7kcFWMylg2EGgkOsQw
dnSUJmv/JNoUBzeasqRqSBVfL9ewPPOmXlK+fFW5q6IPZEb22cRj4WOQCSRwkHPboLYHNNsPhKBq
+n6S8dhHkOWDvB3ZV1wRyHoi/Q2D5OSQu2UnqiNq2DzBwi/+GNI5PUL6XtX3WduBZXax7P+2IyRx
VDazNuo0kQjiHOqmujLKv9ZdOW35DwqvK2kV1nz7OahOPg+RsoH6nI/kul0jdJZiOG7UhEl5Ceu8
rP9QaQ55AtJEz/VgYryxtyAo3EyhYX3lu7QG0+GMo2pKhjvnnsTvkS3lnrQOi21GunbplthEuAqN
VR1CRMUUrlLvJ4oaRA/iGqkkPwFAkYYK9BobJqdJr1vqTTiZmZoR3KcWUmPkSvIQlQiQsoGHxRNO
FhQ8WGs+cQrMYZu091J6VU69Z7ELBg5LYpj3LvqSZ/4v/XSMS2pLsydF1ms4W791B+TSz7zwdNvE
QU7EpsaKAYFfa3cRoAE3UVYhBPRrvldm510YegONMap7/007znvYERGo9fQVbfDiVDBpk+FiqHnC
qq3b+2VUU9TnJsAoDJYfTh4iB+abM3PxQQG6tifYjoiMZBJNG4Om7t7OOayzbR/OhhU8wt0wnLw9
5+LTnnHiuUUhpWjnMoyNJnT80urDuG3Ru4eg6Hgq2qz91LwFgBSyx7fhdN9Yi5qU9hT5t62hNUXr
MPDyB4w3yirhx5aCXlnHvnL4s9fdPEOYrKQ7YVKs9eMm94SupNMbQ1kFurwDfRlGDzu955YJgILa
Op3XJZgenGbshDmIkddOmBf1ZTiT08EeCJ3WzTe2s2THH6th7FLRfUPdlq+aBqv/2R0KVU01zUkG
Cd8YwF9XUeL7VzraURsUC9k+rldLZywIt1X6bD8eIJbFwrOK3apbkjoWduUd7hr9JRXt7o3gjqQg
hMcswF/3AKVmEg6u9Jjo+jVe1mfSb4FhZ5JIvwMXm09/ns5MS4virnmMGx3hbQSdGnSCMjcWDuaU
CP9ok5ixcWqj/AVCqlfNo48QH+JISKg9j8P/t8xhJo+Fr01dmqVl1zmZ39TiEIINBqaZcMjLxtRE
+LmbFdNUk22DesiX1uS4OweW9ITbNQwrVCn/Y1Ss3Nn5si75yke/SYNCEdWGAxvzxuBBNCmmLaHI
sbGy95CndfZ5+yX2bTNoZQaDLEIKazMSqGauWO+EvH9TSljExiP/V18r4K2c2F8Lx/IuxXmtud+B
rtT3l50yMh9FPNnhFTDCRl7Y13Yek94SQtjMEYS9BNncQDpiy9bAIgETaRmkqrENFIO8A+k6vfU3
bMq7qjBU+YRWnkG69BFsCpBeB8avul3Po+qSf+djiM8ZZoyd215BRNVq7hf8Fj3cVm7q0wGEeJT7
RggbPZUaHsg1EMSnVBmCINRFQjGUb0UbfPcjxC6pCa7EtIFrZe7vD/xMBUK3AtA8qg7E7NzIUVtR
WOkhqWV1tRI9DIg0FQuJZtPUAtwSMqU6X7p0kssywNJ/a2KOr6moSFj79dpA90h6Nu10fi83HQ4V
xcf9qKsBDFD8JyK9wjyJezseKUW/gopVDw5lr6AMEVU7pukbBocod3uKopkrcFI7mcvkHwg5Nq08
9YdQwZmJyg2jVKI5Me1cUNvmAQ+0U0kSYJSpOr+ZqYroV7hj56C1iARGu4+FQBLwKE8+IczYNuIk
8xdpOhmTNhMzSy4ZT/ztkWw6KUrcF6D0V7A+bt/psMtMxkid1XCohJq12yOoUy49e57cQkuZ1x08
qF3KHCDHGHYSg/uq4EQMJsQ9HWAQB4ldjggQrb4TcTsBl9J0mWhR2QytISNijC+/VaPAFp0gGEKB
ToHB83D6s1MOF8lEX0j1Ov8+U3DW/pAM4j8IRgNDfhpz17xPISXRBB9q6XGJ3iVp9vcAEOsA2KGx
Yd6BWpttXow43ZDEaR3S9MCyD7vniG+STA6AFKYHSvcUpvESRiWa7Uh3HQNbLgbYk0Zd/3W8BMEl
0m4B946enu8/hvfD/lTWNs6tni8lLt6Bct9Q3EvBeI0jiAvwS6rEAV9mLaMZKBwO6tpJRpcvpJPY
cZDfiGg7LwCf3PaJF3YQPfYEVGKwO1RPVRxiAlRZWciwOVk8Pxq5qjF8DrQxMCnG9bhIEMyFb6j+
r9J2bg0wnAPaUGpOIcMPHKPsqypog28nNa4pFLcy9Xw22cToGNv7Qr5c1QE+kqBGjMrh6TGKuHgM
1AkPwLEH7g67lRI+GbVTWnkKYtpVhhk67kD0UABZeiD9AzjjzrL5B6buZuYXkSnZjfD6JjGyjcJ0
vfMEdMfR9/L4Fp7MmOIScv3YGEUr8WQfNnQLD8KgCCpf/v5Lkki2qsuyWoFY/UWzJki/j+wDtDPg
w1YLG5X1KVZqkkR/3da0hZRvaEEc+wsD+h9ZPhnM2C3rFx3ZrPmI0qoLFQxA4jUD+L8l0z0Dkryn
QmdqFd4NolnpDMjwpU8jv3cqmZFkQZnB1Z9275aLy7RyTyPdfAHz/+6eJzYfYnf1xC+kZ+9rW0BI
vg+UdLo51sGByAk7G8jcd8WBeLuacpHswqDAaZb5NWJo6N6dUEsTgRmBkGTaygXu51aal4gR0meo
JHD5T6JMuDKRh17AmdIOgeoSrZP9TOMq0Vqv9/F22xNjZ+imEY30ibaplBjD8dlGoF+JdTYmXKNr
Lv9q/nikFoOD1LzSyZkavhEUM7PWGw+5LeBgHW5tBY472b29FV7IlpWqwdy8Beew5RSYc+lSojcy
ujBWsWLE94tesQ8d1yXsPUg+oeIKrSwEddGjSIAizc1EeKfznBEyiR+A6x6PDirrc5v1xm5Lzf1/
dYUeUYjdv4kxFiHvKKlEM4eEykEnIeFDsJ3wKZYGISOWTInSHOpP2/Oe3dCBLtPbP3KK37l4wa+r
D3zamS/qQhfhZ3KuaX8Ds/OtBQsBp71WM/CtarEPCMhNpkI4MD8tUJXfOtHv7N7/EA7/FVBhBYBT
msFRxlVVOstKM+t5KNuSgWUrA06RQUM0pALdje/vauf4Na1WscNLxyu2HY4lm3Z270ahJxiRvcig
KmX153B3KLz0iKgPSQdjS3v0yds144o7TcsctG6i3+BAPRTuglQgD0Jj3fnaJpWR4h6cYGeI86MT
u22yLL6Djf6lhTnJfcLUtSJGl6h5KsVHfSmgbd03vtWl7v9R/juw2iKFtI/qcMlbpImcBObTbU4c
HZ6smy58klQMl1a3Sdzx3aMryaJwIdzFOr8Ysx6TcfYzWhI7UyjDZAJFfrstvzunyGn0dyQ2s1Hg
eRhgKRA2K5+Tvuqy4YSCxaQCwDaW8NEDYJYm0E/FluI0J5DWqO9fQEafMh0UotS97ylqfYZ0vSR5
BQjSW9oI6TECpUeIrb9P06QvVa64YtMHeBYSr0eJC5aXILUdoysEtOrNzL+JqLB7mYAEygISkZVt
/zTw3bzGhqX0eqhQGetbIBxP5EisRIHjTPBG0ol0LeGprBkBQBxxf4ZYNQxU4qQEvWAavQV+qVdx
Y0WvZ93CCK9a/rLeC40/dpr5Wy7kAOcbmoeftlD60UyOZ/fJK3O6uEaKODHr/7nOMAdzHeyLwJNp
UwpAW4PLjg1whW5HyNypRIJy9myadnspI1J/KE6uCrkh8h9vT9HhOqrDOmxE9mgyGmAbtvXvEN/N
AWFWWwVFMNVQ9aWZXFKVJxhpkYdeY5ZJWWS+64Iy9oZVPiVjpk2s/HUUoWFGeX/oAwt0t2F0nynM
pHl+jsVhhtUqBgvSAzHqFuI7lCY5Ai7wNARyu4Z7ZXRvSw3ewGCk9AAJH2dBpDOOeFb9R3HOyCG6
whusvbAlUkl2c7xLhQtFIWV2i3d/AoAfqADFEm/dv1x192Nfh7dFp4ZWVN095vDol5m15Fmgp1MQ
j/laSk1ALXkj8Up8IqP25meXYOOa9teA7//SnUd1fu2YIiTyXemyXOnoVfMXj2sZ2hYDPGCaIwtR
gVsHIxdknThon6LBIDarUEIeMOErSWqPCdK+v1lxId4Noc5XplojKlHSHE+o0Ia0tEJu/KfkU03k
dtl4FGS6FxnHbr0Qk19kuLXPhoRYgX6oZhgzKwqIomlbFCafPY5sS6miCr+HlargfVCOM5WcCIEq
3+fawdbHHHrUvqQJJzCWbSlvPzBlUnsiWrRgyLS8qs5XJdjFykzEn/vceLz/xxlvCfQtFrCfnq53
rpl4ytyzLsoR5bJMNJzAN9Ex5yYouEsndhaOk33QBc63U0ietTuXZ85MU35LPNqA6frP9e7rJvoE
RRCHEJfg+KvUl6d5g8+gTuFkfoRCmkh6Rh1cJk6N4f6/8jcec0j0TmpmS7Xx8TFFYWhKpRF5nyXZ
H63K6DsHgD+QcIDFa6EuDh8/LQPhSsTWdnOp3LbBX8xLnilJrZ5Tg3Ac+ALVzFD2lpCEwxHMohBx
Mgcw9zpA1/oiqZpbyG255ZPMx5r7RpYchmMLboumYMKRCHHZ9SNFtZuK/dhzN4uNAkkT5UN4Psy9
/fd6TDCqpGOMaz7khbEozaFMQoLpBs4jfvxF1PKJYZ19jUUPrCnWmso4tKY+6MciapLkSZ5TrA4N
qft1seYgryV7bLg87sANR58w3X3nztMvdTxArMfwgwXM+lVufKp6YVt4XPWz3yOxUlq9XOYq347+
bNIek+vmBN20cbgGE3abQ2vKzLIS9ahG5UxOOYfP8SKqoP+X0yXx16aHxBHeO/BybnXWQU73LOtB
KkO+TAnug52lOa157YcTBf0NgKFJRtn319GrDroZQWR5AM4BSyEUMe92wa7rlHjg56fSQ78DfBNJ
03qV9VLglqtA52u5DF4aW/yTQNN4vwHFneVcB5/CDNDpzTybWh1qfPhgzqJz+jr//R1QZTYnRs/w
Z0ZhoWkOU3JaQCawSR1KskKS9RYa0rkImPELHSqmiw4ieLI+Vuye2hKNT6uC0RKDbNxqLdkNNYER
U61q8bleFaimSbbACDqieqImKoyaDS4BQuBlTrChdIutLul7lvj27lbtOdsqW1IxMYdpdlCHp9wl
MyNz5Uw+PveftkgRa4hJ52Zu5xjrAywspnepu1ZOZOnFYRAk3dsHI+MSBCtN86RPcylNm+1KT0jf
c8yijcJ6Si1V7Qr1L2MLNAkYcIkLSxpoieGuJ2COo5fPI3Q66OVbUAOoblbm8eB37DQoyMfGt+B1
RrwaIc5aGLF6zBDRG0ZTk95w4B5BhJXHuNIKHWHQTtSvhJxf0nNwg0FBV+7Oxtzu3HabN33FSa1J
2qiGLearYZHSAgpT5+5Zk8cFUTFAKtgm5RLYDYhHvqODl0lw0ITd2YLtzeF4Hy/coefSa3RmsrNJ
WVynR/y8AxBNYp9hklTyUQKjnXHHfXqi/PKpiSAe16Y79D++ZAYsCeZjazHS7nT76puVAlwB72LY
8SAbJLsAi+2ihsUiovNN7zyJl/v9Xa6xLmt9XKLo1JE2BBYUNqew8VJz8IL2Q4uLNBfAwgx/uStw
/4pAIZSw5t2X2U97tQllIcERrnoChpz8yHZzP4lAqFP368yZnWSSAUfDVJRvfg7dd6cHEw808h8Y
hqKeKXqJwbbHm9ch2+YLnpKouuv9uF2UHeVC0HzrUgJU9Cxz4t5jtKn/0JSGRikq4Z+pFyAU/EyU
fqqM1tSxVW39RH89G56BFaTFDRCkn8U5AfoMrkPRymhbO8b3LRdtrzlHlrBJ43kJUXk5fO+5Zed9
7urwy0dUBroUUGIoXi61HKZtcRJ/5lr+IJ/CSq4fBGsTIcAKLxrv2PDtqoUmgZXb2xoIdXWpuSOH
DwVHZuJmHAjfEb1SDwaDqwA/0sMMirDGxA5+tTtZoz+Ds568dVC2eR57xrkwZZd5GpcXgOZwjih6
B2p0P24hzueBw6ZT9svSPjE1vEjZLWYiC3rHXVyX5xmktbeKD9e45BF9ISBtBxTev4A+avih1TEs
qY3zTexHMf9WwbKC+CUS0N+hfhSsGfst5pU4EfgbXnuUsrn6sxQYNEKDj6d2mH6bjqt9UU+t3ZJk
2YIQimBGI1kyhVwMo+/MLkIYBt3JVpCALuv7rfQs/TdsXDWRWTE5FUkxWl+pswN75kCiCLCANgc2
nKWqf69OwgKk8UD0y5JCcbjbxMmyqk9TVdvSXFL7p0kmz0hP+8bGhD7LqbYmDaGoo5AUpHMt6y7B
zAHBuhW/TRAtjz03jOG6KqBYovH8xKlJQoc4I1Zx+3ti0tohkri9FatuvTGKLh1mF56YOM5dgP/P
mV5zNG5RM6CjaEsDbNmY1uY2j8hNVq6SB0F1uZFlQOVwfdLtgjZ+Fe5d2XPyHO3ldB/cxfe5fBrm
7dRwQ9bxGqzlmlrFV2hj/iWu3t8KMXSV98lh8lfArjNOJSGEw09bYR2AHfqv/W5SAKceKpKf1fBw
/fMyFAtqfbZgi7PtqO+mdivg7jwqbDSCcBsol+OddWoNIjXHHsiyfvhW7DGNKQ571NnIWBrDTJiu
/17waY6sodbLZw7kwQdq9tNYOOiTMgRNTvcBeQJodfbsoEnKYQpPB5noLhNF76u91KqpDMJM9Fky
E3znGj2dWz32ZHaYq+JdcIkbAdnA81UeJb1+K2K0OiEBJY13Wp4Dt5b6qYvKDeQNWF1w0bcRezRe
SPQcQnY+kiBlZb5gI91anycuTzF8xYvW+HKWDnZFvhOyE/btB5yBvFt+lw7EMa9kvIO5PsTQBrPz
mNChIg0TqBsQf0IADaYkJo47laEjpY9hMMKAHPlXKDvwNv1z/wtUGpYhnR2Dr7va/CaUPcgjpz8o
QnQqA5L2gDZQmYk23MjnC/sTkyh+HyVHRIjoQcQs6fWUaRmY/hBMAFmXNWeWTb+D04dgD+ov9YPU
kZbKjFQVHF+WOtWprupEc27MVm8+UGGNuCI9EXeD11a+ZHBzZTlSv14us/yYs1kcHSIlEMJP1JLh
JmGlq/QWvuwBCiNvRGf4WEwJpN4/akzOvGYstoBsLpUldFuUKH20tqSAAhoNoJi56Jh+HPFRAT7k
r3iRgdPNgFnaLDUN9+v573JXwUaAa0b8U+3TqaDH28vLbA7Kpdmal8Bmb9YvV3BL7/J0TJeJu894
k1na96gX1K90rQdQLGkPq/eDH/45g0Nn4sFucLFbKRH/yaC5gboedca1o81ccGfZk+QHne2STPpt
6T5CiQ8WRKRuHqsyMI0wskxtAolwhBn54wQHcJU+8h5HQK2Y5nvzh1nRQK6n4HENWH0lRp0rWoTO
ufHSFKpEV72LweCMUfzcJ8UV2aKC+pWhdYVnqPS1OftJ8Jr72m377Trr5JtIAuDkK7UIaN0lBJdo
/wlQJdlBlps0daQwEt5ytAYa4yhqx1ceZ496rBbk/KkDSDaJMfKN6y3xF1+DadUZ4oN23TCdg9F8
i8RaWm1NQMD4W2gmO43RpbpjRxKCWkOxtu77OG+4kMDb/ZOHTCsY0T7OikwtbOwSsf8puCBWujwa
jPH5+M8HZTVDtzirpaM93iV8lSpGKx4VhVlAp/PLWNjjCmW0rWPbUEux3eo360aO+qeIMCYZj74F
PEUTbqopk7eZeWBXa9usOnqqTp4H/4lSNQZHvNkQQ//v6i5enTNUQZr8jFTuLUnfBW+M9D395NYi
Jebj/CpeFxfI6FGEJMYv2mAUq8wq8lfn+KcupSMab8juA5L+Iq/DlrxXf7aUaNZM1Mr1L7n6yXEY
+V7h0D579ntVrVOU6zJefLNkZaom8rhVnUkGmkyC+jEZsAjWQWvF0V9SecZEcke4SMzNDqEvcooV
UbKmXpAtnoIhRjZ+1ARboriv8gPtvp/yvwDSKpcjLJ8Jt/Jlf6EXINOLY7GmzlG0kxkMfGF3EM2Q
32/oSfZQ+eCXWCAw/Yp2jWUeis/rsde2h06lhZIF2YmTCDVD5doZgT/EG9yObrgnBXoxNW6DPZCb
htVzKIdUDp+xJL4P/bBjPUlAccaJKDWsNNtWrNPghbT/L3fXgNYWtGQXXF+q25BAaKZZLkGeZD23
jssgU32E2ctDBTxokouRrdRZD1VyauS4ZS9hU/o5jXX5Y7cseBCTkPfJQuG8cnQzTTzC84hO0e0h
K8ZfBSRR95Qx4ikPvDwXPaw7u9E1A07+ByLdZAW2CpEICfaBW/XQLwp+6pAEfTv8L4r16/ngRbkY
U1NZX6i2hH++KrUsb5R680Pcz0YrIyFnQhw2S4JwADEK+/DKNI2B/S92kvyA8bqDbXx7ha+SfEwp
g9yGNyzkSPwXgyMRV8Cqx9/dCu1WYmcrdoNsRXUIgalNEIprRcBIOeSXdR1Vh0MWKif30kH/CQKX
J9pUwC4yt/t/HKYaBZKPcs9CEL3IAykGF6Soa4DkRQj6YG7iRoCh4ADY2kfxQwHthfcuZAfcDTqI
Fl9bCtf8SXYRUZV/nUSibPfRjdqoxnuo0Sr8IsXqLRHL+jvfvDC6c032Axy89rZxYCugUoBfhhy4
N8aKGG7GcRJQx8dQaaTjUQPqKXQ7N43uMS49sCf8QLksEksDfgllT8HSaEg5LlK1keP08BESgoRi
R5DayV0ibxicLrJg2zK5D43erfFhmTDmBCgzSPm1dnLWxhIwth8WIS5gnSxI4QTsRguLqcb3LL+g
429W21oUDrsJsSGXybPWVNgHteXiTD5COUlghS5ZjKF1CGysjZlrpLsJz0MJqmm4M1b8GdZDhArv
JiAWGGRVy5T2b/9yojpR6Cbphs4cTSX2DTftcdFTL9AZrzrbNOnhcqfBjn4bCpaCTLzytypCsi7e
bkQhouwSV1eMi5+Ue8p51TCFFQcpRVSeAO+eHG0PZd43wnJnjOHGVSYMz3hR7sdmKJ+4SUKzRmDA
e1iNz031mI/aWWbFOtcnG85/vvrnUVFX5GYIUDcVKQMA6sMoQnYlXw79JujdA9vzqNQov5AQIhKY
AclWbgXXELDJ+8x41FRuLneYhs5lyA/jlvZhtL9eVT1TnxIzyy51Fby+G4JaeLKaVRNeHWA6PqSF
0aY3GRtACY9V0GLGssMjogIVVyi1PItd2FopV8Ou1U8L5bCR98HobvOWFHdf77Ea8ReG/avghzFC
S6FOsRJlDRrUcx4JS6l3KjAypCcaM0Qp80CzJtVGkWM6uHlGrCWg5nA4n1KGMJAodMgxHnU6ww8D
136Su0mSvrLbFgj7iMuw1SAlEFKd1B9PzY3gS6ZM0cnbNVJcM0X/lGPYBuRyR4N17/Ey0C5zoND1
8NLZ5ZhUukOwd/WAdf+8J+WZ1RT8/0WqTGwo916Q7+U7sz4ihWv+2MH+lU5bhAx93AakYgYJ8m93
Y0utlUs4Ut+C/BEuY9IMZ818fODjvaRYbucf8njW/9JvU6EgzjQYwzV+4TDXgkgPPn0QPhdTyoJ/
exKD7K6NJNeIMsXr/hCPmjz3zakcqYwLvjMgOip9q77e9FrWczJjyhb8HGFDbA3lEYHt4TJxF6O1
SfJcshS31RwJrppw0bdpHgdNTJo00yx6toQnkrj72Nlb9mI0QDzl/lggq8h5SFHBHcVx/nmHgJfc
rQ905PIJQpHgu4W0GstUikyj3Uat1VM4KcpuMK85ViB1w67JQ/GDeUjwgNF+glPUY5M8Ns8tRpR7
88QnPW9+r9E2rm33jAWNaLNhFY/SkLvPjkrD5WJ6jJCPFmIshTOurP/t6BePiS2/wEYM9PpduDr6
K4RAYmZhSMPqQgP4NOUCBykaPu7+7YcCGIIg6s4CtlmQjIM4c+8Aco5/naYuumtaHkxB5wRc2jiK
b34JYdDAglhWkc4YJ/UUWVGe33Cc1RggrI37nYorZucRdiRT/HlsxLdoRT3rlbLLSTKEpTmZWHp9
5ql+O8C7AvbgvgJh+dOkS1U1mYHYpQ4wuIHi/tJaf8mXiOr5Vjfp7w06FH7hTq8r+E/p19Lok67U
hQD30st4thGStiRmqwUC1Ch4dn7MWQa55PjAudLQU487V3ckm9T55okg8oVYpJt7fep42JLQvzia
3EMlz/XfCCSaCAcaHkN79N+deQRj2e0HEMdMkCt0WNcMzHKS4qumCoAnlgGXDlD5GllNKksfHERo
tWRSxfSTKBtqQtURGegm540v8DuBiniq4nK3oUiOIfBfcF7WSILArXrzbhUG84vDi0pVuohkXTLT
Us1pzAcKR5mKCxZvD9jdN4KrdKk20TAwQsniMI8tZwM3dBPTsoffnkmgbNepBREP/R3xxiaNLyty
R94Ims0vwi6EhipI5hHFPJLHQCLuUHLPkNBPU+hv7JVBRe9h1u9XnE9j7sdp8nCMA5ey92I+REBH
rMg5RI9eDJHTQkvwARPc2dm0KFJH10c2XxAij0ug5GimVOZxNxQfK+boapOv4RAwrK0hw93LdWC/
Ifr9RKy+nk3f456ChscaPwkBj983mDjRxH8zaIefjXkyIQJCbf9SEOtKY4PtEVrAlf7lZDnu44EG
VFpS9iFnZy17jgZmPnT+7BwA5/cMO+sXd+aJnsqo5dkhr5DH6TF+/iu3kEB6RrUu19KDbSnbKLIi
uaIJn2cEdVBwe2LWu0C1gEETQjO+El7fSQmBINTWogohOAbqrg7vJiNMPERnW0yaDPEJdzWwAk2Z
cd7GjBGIB4d1DgOEyuk35ztPKvhN98Zb/TWJp6Xkh009pUU2SGOXHy5InHL4XHx+lMUFeLV/ucns
kC1dVsuN1htyioXdyAeCK9jF2uuVip7Drhr1UapSorHwed/5nnRNUPVg6LogAyfNwMvujaykRMl2
Zk36HGW9KoGOY5K3OW3c3AOAtKXOVn8omBnOCNjYEHgv78wrttM9KXJ4eRcz4qXrL90z7JtmZB6H
fiFO1A0Tg9qP3KEzaGHHtK5Ilenzztfne+SvtPTK+h0/7J/f0yqxKtN9P7QHpCDrdDVOrZLee4/4
RNFKHXEyX+svLgBSotGu9IVkdQ+RtD1NUNex/GKhFGHvf38VPorIf7629KnWq/i6DjJsqLbgbcwz
oDY1Ic/neH7qssSxGXDH8kEdBruJhpQKuWvlh+fqf/xcdl2p+RFsqWm4s0R3+UgR1uH8TJIe1oRm
vCAjBnRTA+2GW/yXfl6f494rcI8ET/mlZ23uybGTan3L5vrkYzjdlf0Jh3ftA7R2Gz3ZCBlAVlvz
OxxOnANRKjfKQkwM3KCG2CIIRbu9dnMnGV+wRTmLeIFaaj9p/oRnIaGFnq5wBBoSpp3EMtd1QQrA
VhCUHjXlpNYTFvwGbeQb/K0fLy/lYtm15CO3tsjbRdCzmSUXKAGyuxP7O8c6T7Cp5JhRvKy8JDwH
k/WVjkStpVqY7/l1eMpSido6Y3I/nUFM4OS9ShHU/w+194zj4gYAUzIEH7TJmBDgJ/sTU0TcI44M
0lvfmqQTm0EL0TSyKXPt/CC3gDBLBwVxOkStQhhLHGBQw5JPf28810NZ53Qfnn6u17IJhVh/SPQW
AP3YudyQtbdZ4cjTqz2AsqCbfnCrecB1Bo8vMDJb2nZgxgist0ymeMcapPFnP9MtDk4dhy0H/awV
aHC61OJQcP7Y2m7mN4T6+xZaQlFbR441wS7z1MH9vGP9b/tfPxdB81E0s8Ne1jSX35Ez/IpQl6Jl
jQQhnAD6NajjBMeWaizXtiTxWtmBH7PHyQOKE0qu2fTASRPYmCcB53l6vHjcR/4V5hMzpp6twhwG
qFLCIll0vQk9eMSU+aIAkCjI+06wJlGOhswV31lgiktQ/iMng8K9ulmHmWrOcB+M+o+gPbi+mQMU
UB8lFQ/wNhCqw0JGOxCKIhxWSdwVxC805oUVn/iSmntmUXyU1zulK1/zyV905Nhbf+PTmSCtHj/D
VcV+r7zdIyn+Mvm3sJOjihgtxUVrQUjEqx4agbKJ0198BfUsLQAAUj2tlXXkcRVIzJfBMR6auN3+
yZCD5OM3vYHdefBApeVgG/qBvO2oKlyiN39d/Vt4tGKDFCERjznHhkxA+lqx7z1j4jqSiq5E1qx1
eMMlKQltcTw4cXVe+OP9S4/Q94/6WU/RffcTKwscsGwj0gszjq6xB2MrdtEnyy9lDFuI7DZxXMxA
xucwhi23+apQEVzX+tZw2+ZHZ2i1pCb5doBt9iaWtFzOz2b59OK2KfoNUrvnHLmSobmUDIekOv13
KjkXWKqWmOB9iOI1qFG53Uf3J9kQ/4mr7gL2XY/6p80KVXooXgUcg4dGi838PqlcJ3QB9hB+mODJ
M2NyfFFM2pnbwVscq0C5OBIdhDlG/cFAMb3khkpy0fgDF0K+iIEhoa7j7QYMw9YFqG6AH20s3pQ9
NOAZM/UnUs60jYzt25/R8dYrzozsiE2P0zeiu6gNnh5q4uOFrMTqNGVgM1M+Ls3rnUHwbTNYbEhH
15iRpdYedpi+Ex3wiquD0ZMV3kaAo2+orXnfufz+ySPWK+WF7AugC5fFR87AnM1TZOEQOpuLZkF3
DJvzPQNASvnqIJVcxZnIkEThFYC3YDP/+X/Cis0LPnqBzWZZppesLeFV1xp0llir74CDwuvfr6jv
mwwxw31oUxJNbpLt2b70H2gR3Acq5kat3ffjE3Oev6e6a3exMTT6l6679a1q8Ufz2otYlfrFs+Vb
Dyo6pH6nIZTvqyQ6JSaRoEpttuhUY4iVxVPZdckG2iELYTRd8z3oVr64uSyEPEBVQEgXZfrTTRbQ
VsgS0ffGFheBhaCQb8yY71CH/MN/NI0QY7SO4kVWJ7VX0OGrDCJ03Ec3++NH32jLsxnLG4dlM/Bd
ru507pvHKa1nzPwN9koY2+Czn7+H0zjQsfPPN6VWOyiX8Q7/CqJnk5c9UYWfRUHg591i+sucxfii
Qeo7b4oLrp0jmFcAJsV3xo1HldNemSUo/3a5lNr1hCprDy7X+bOcNUmlHsdtfl7jdOpzYEEX3rjE
uTD3kOf9IpJUL8TLne72sqoz6TcM1HFTy5inHBjivhkcWl5t1lSHXm+bfjCEXTVaRf9fYm8Trxys
VtSpajg4h0a7XB8bOPWYsWXaKiV5F5iJ3ZMTzMFWWOBt6pFy2pw6TbzmMVUJTRHl3NEsgNWJ9d+a
e6nN/ElPeKOvVvYkV9GbiaZbqZ6LwCkNvOCQYgwYYdkwe4EmAD/2QoypzGk022KJph9P8+NTVLfX
vvsBxhOmj4DpRTIxZjRGgcdu+5aFr1uG0JtXGQ7V0K04VwXDIYIdxI+hPp6Bay6UZJ9FcX2q5/Jn
ZshltTb1OJNtXjnc9jGQvQBmmSpQUdK44tj7iFpMZOvl8SJe5EVKL9uCpWFQ9wtkhn9HksOmoSLY
Vp2j64sttNUlTxlkw/j20HK/0VNZoVdKVEu9vj/BKvgdFBadWnFnOt5U0QfHmElHgmN/pRZW7Cbs
BAy6jw9o/Fp7UNOTRAKlN8kAdoc9KaDzKAgZ7qnMkTkQH1J5LDpE3Yp2sT/ZBWzpl9ErxkwVzSk/
8FZYlHIMhDIseRYS5OrMp9uAqZQPP7senRy5iIrPGnaD9H6m5ijpwqpU0YTEAbBeeODiuaNdzT3T
78Y7dz7J2YaRa/UpF00ukRnA+xUnilJI9Zs/HjmZodoiGkazMFo6yaL1qGnAbxJmQ4lfZh990ULQ
e6bzzcySIupRyzL5I0Z9C29B8aWvRmVXfeRlGL7PbCZj4d8yduewci4WS65Lt3HZst6VYFEXYZUR
HrhrmQlgEkvrhcVZRdyR/6R6fKtu6O/u/xdAbdwwCkZKHN+d+mSmQEJij/u+Y+wC8rKtD8z+HuA9
T8ZW5Qk2IUAfw+56RvOh0E+9e5y3hVO5RolR3a2e5L88y7bo6tv3FLzgL1dB5hv8MlxP+zDpVv27
KOhQn/m7ilypsPiYVB7k4PdLP8bgVt9dsZc/QL96FngUn4siRYAnfb/SoJTLmgOKTEP2Ugc+TT/e
iKjmH0HSnidrRiYP3CQU+Y+apDdsmeuOD+AEe4yXoGakiBarfA93lrmKUmhTLGkxVEyzxt0PJw0/
rK6JGyvO7nEo9XoGP2S0nBY6gL0AjKQEtcL8SIBwI/lV3GkYI5NoCW2+UaI0VGHETZXAYbYzgsUZ
f++KjzIm8PmjPFuNNOFfl1c09ucQ+7I437QTFpD05ne54gSP3daD5J9wwt7sWaqC9fuF65CdebCz
8BVrCFcT5ucgbPhXpuUhq2X5oN/tsV7idOD7TdQVRSjFIg3h8cnYtS9i7ygqBh3+Y5KKxkrLkmes
xDZI827iYdIdRPlkIy/MzjkLZTwiRnU5dSjHVzlcykYPykiDf7TaI+0/zJVLR3G6ocRNUFQTgYWy
uVf2J1JNXp7DQKmuscOO3cuI4n+qhqq09KY6UlBnSjItwDOm/q5Yoi5Ql5c57tzrKty67ZES5MaQ
UhS/pHmSz2OQpjNY+oZ5fozxkDsi0h9U7Fwycrk7FfuNf4d9gIOai2G3sjxI+gy3l+GDyBuF19z8
dc1xVys4IBq8XL3orX58lp1QINb9DkVMIVW9Xkzf/FBZtcbtQtfU8eP751cs7mfAWnU67VgJx+Tr
zilgzANXVkWbMKaTgGeby1j5bkSQBcO3XgdD+1V9ITb3ZLbRSxp19xAC/kDykvrixLnygELLi6Ob
gJnYZ1XH+m5QwC5p8AHGaiBhNyrLzit71wtYRACJogwb2IZy7P/C/qsalGp+ifVR+MgymiMOqQBm
iPRdvZce1GLRB8JC22/xm13IpllG6+f4ZKbr3UAqVTlNHgaRcTqx3JLdt/suClJMUDHPI8SzjwS7
s5YwOJZk37MkpAyJUHGRe8gjbxebl498Dxcd3268xjxnwin9cdVl+MVIGi3sod/dG0k3qnUPqIdj
PPpcMq7Gr8rj9xCW5bTxdvu+KQ0bYWXTHkF6xdeCorBd72DuMo9TUE4hbnNAUYoFj4uXVvDwEuQj
Fy4MMEk2NTHy+pmECzYthHOnu60rsSUweMeOu3z2X5A/5acPT0pSD+vqAlt7En7NRBbe9or80QIv
YRTJmi+lvlBnt/BqlxHxqcy/pPGGsldnQK/zepRk6yHeEL4QGY1IzhMhMQzZoW92CE7euhizAF28
Ych/+ZFOmK0TjHPj0JOsAv8v0hT7DZe2E0xZmqc7El9Q9WctkowRi0U/Nw0QmcTpJNNuGhgXD3cH
HSbaW09xemssHG85ZfIuBTbu8glOi02L3MN5XObviyQfdYXsoM8uhtHBvGTKofmxCz5C55jWlomp
V/w6BA6dUOEKQS2f+njf2nRGPy+0K3clo8ber//1CcrDEF3ZfyTt7RMPb/qhpUe2tUikwnnLZ3dZ
eSmDiKOt1FA/Pdab1dlNk1YmIYLD7rg8DOJxO7sIQsD8J+I5lLmDBN+TRJi/CPfOLDLmpV187KWe
YoGncgb8Y+4KZGZpLP+fimSICjwAvjDcXxGAHm4pRWfNeAhMKD/MXdLqX2xBORTDDr6LPUIwY2rX
TnEXjHQi150AYVtUy7G2LNiVRHDdteeLXy2gw3MysMV8+DUxtG58ClOW8MddXCn+Y3HSU75O7AN5
eLUOUaHDOSzJI3K/hl9R40FIAwrcMya/c1mluno0mOJAuv+n5V8PmdkAR/+UjR2J8MWMtHBGlNcd
7adzZAbbdbbVB6Q9GzETGfU+51xkPY8DzFViG1whzmscMvuHYsJeDY7CHWZLs7q3+4fpUDwgw5DD
m+kTTEjcAzJfKYytj3wHBaX3tlGqFK7gHXCDKkxQVE3MW2mYcwcd43xwylu5tX3Y724Kfo+ckkWZ
jWJj1TloBuVWVxNFT+CsTgkpPzgl26xbbArmqHjpkFITICwAjd3otZ86e1eCJDsw07DSzEQihX1l
GKZMjyHG7v9kqNBbIRBTlnmfv4xBj4Pof9XzihOnztEMDNgsNMrmACcc7GtitkkMm/N7pcxLe/9U
pI/OmJN1Bvh+GmKG5ZlGckDmBE7F7kIi4bkf0KQaPB8coUL8IeVkxu8j43RCO08b9+7cZOQKO0tD
5M6tM8zb/Ft1jdioiA6168cr8aZSfe+lOVDDecS5NRLC1+ILGzZbI6bZpT0xCaq0Th6dU28Fkoqm
vi/kJg7C5TJNbGvGBY6z7P71Y9HhfYdTGLCU7GO1L2WIKGSilgll+dJSaJHhqwhiaZzgGTvNCmvk
G8/HpP1lQFD7Qyd33JPlOoFu+RKuoYBGBPqQoci3+EHD41URZZ/UUki+5at5HgKfeFp/eFZZBJxy
njcyMxalSqkgebcQdhc7pF46H1Qj6tMsKlnhzhZl3tINJ7VJJFROIq8TnnBPkyCFpO8rfBEQoiqr
S6EDpwpOV8/jSUJZrd9J02WXGt5hKRiCuBngAkAFxEdqzNUJAUVlbKP8ICyPO1AzSVsWiCJITgOr
wVxUrI7J2RhFKPYBCZz+OTHL8JRp3gYtw9KBX36Xg3wsOIvTpPHdujOP5Gat5PCfiI33qp0Rxni+
wjroB8AixqsW86QzhsrPFbqsfV3oDlZ7u5ERbayLjvfIo27ZgEhwcaCcBGcCm1hnMn8NYH82QCK2
EYvXmYA7MrQaglLmxye2cUHfLadq0NIuYODUuNxRq5NNiAAjh35UaxpF2x9N1fWDNzsP8eIB3rHp
3w6CYghbJlx+HLwqzCjKdjKICS71ZrX7YQ32ShBH6o+2TFmCJbDGJHKNVohZkMWlmkNp4ULQa5dt
azr2FdEz1te8T897lWankZs6O6/w+YyGQlOdNEBAJZk5+lwE7OJpJYEt2O9PWHCmO8AzfUzlohMZ
Y6oImKg2paZZLxSU3oAG2cEE2kftq4CDwu8urYZvRmraHabvTiJFqGRZoXDE4JC+XTRDE07pEAjb
3s0cQ7VepV+ahgRxpqT+VUOEERp/pbarTl1W0ChNIc5vNB1UqNapaig5XkZLtSRrRWKVmgHncFic
1ywlSWM0373eA8fBCzAIpi5YjxnZjbGIJcZU2feNEc14kQhGgyWnxd9COc7icRwaXjylGaaSJOpc
DY7mjDnGbUNJ2Xwr2TQZtHpdg4wj2btFnHY5eNQuMn8DG5hsKdzTIxPCsi1aS/TE55vsBVfCX668
rsk6CVmiEp9Jpy5UILIW7+apFw9LFYrxpPecTpbX97zIOffqou4lUchEp6nUbwvrvkXSB3/gXCx7
36Eo0FcqbQ9Dct6axmFWTcDrL79UcKSfNE3nMAlxyMdO+UyJMPPgVdBQRhcb5/dzipJO/DoESvKt
wicbFxIEJqASNljeoUXzrjKQBujLBtulg7EFxBZZ2mBlv+vmuJEX6XqZee56H0ZhtPU+NhGNpd0g
b/uRfbgUMvnY/ob54kf4c+08qxdJtUa21Z+7qZIGdmZI5O7T7AHvfm+Ia153WPdmaNqP/ca4HrOQ
A/xTviWZ4OTxdq3jCdVpRuCFCQ566lFAt0Rc5fmvvV/HzMrE2B4M5IkKzaDzOaxYjfeS9Ya4YqqG
ewcEWezpI9+7WlrXXxHEN5v3HLDBy3Mn3/2puydCNY2JZQkKZK5fbP+aAmIBa41pP5xdyZRrZnjR
hLyICebBcVhFlTK5rcaD3UXVvXJKRRBTzeJljClbshKheEh0xB0YuZrpFugz+b109PnvylXZtBIc
jwqL4gyeyyhzpg7pEHlLQmrK9TymK2EoR23qV7AgQpAlVek6Jir2qKaPH9cD6IG2NAYP4KTIrV52
83//GX9zU+y5zfOtEvsMV2yllNuEAePBgB8HbdeBWsw6N2ZXZuCaK+sPwFIvJOqSvlDZcsVOURcz
hLGJeNcleOrMJDHmfIMtobP7krvhEQYNfazBKHr7kuVZUT/53JAGNiiN9crzMdMyDQtuMQZ9Pkzs
tCDHvkst7lmscDUbtaFnmdsAEL22xl3imSgffAPPvU/zD7sp1XWHZo2bGlQF/9bKHACmWx6oApsp
DjnFSTZjc5a3JdnnQaDYoR7127wHMWv47j1ECB0jWVxrOC0H+QdxHvqGPqWMji1mL1gl+FgukzTs
gMXG1bB6SWKs23XXhNTDOVlDItVlabi0jszcq3g0KIDDYFar17n8DZD0muQ/qYSLVd1WjVoidP+1
tZNmAKA3zhQS7VkufVjxs/CkQXU3mBgQ5Icv5kuiRQIetyFE83cVYCGXzyldoASdd/IpK7OP8lf2
U0KQZbW+YSMhRrikihT1J6D87sekCDq/h10UkgrVZARsZ90tQHcjOLwadROXaEkRBLzQZ/5aKvsS
tNdXUqcGcWLvf4Ih/Q0gwEJ/hzVNi9WDr/D3deFBg9E3YKR5xkpFhCOCQiGDlR00ZSNPkurDoKZ8
w9gLwQ4Y9OvJqJT8rsJwf1ZTURY+YDtZ8DMAftJD6UmATktDUmwGjLYJhFt7PAwZSREadvntdsGx
r4U8PMPo7u3pZQdqtPC4EusnT/nfJoEEVJ7hq9yfpBitZ2V3mWiHrQ+iQj4OQJVjE/moCxyKShgH
Q++kB/Qx9snNNkEu4Pi1RZ6OCgq7rmdZYd2A5ZVIk8SH34jOmHGY7/8v5NMvAH6fxRnOQKKPIafh
2UncCWXn4aiUF5YX5XFO0np/pT+7qaxK4frttoXlT2z1EzEKIjskq+G8V9cAFLcHGQoTtCX8b6BM
z50TK2O2b0ARQXv3QOQa02/CKYV2TpcvhREc5bg7E2iqbOm5S2MCy7E0KQIc7n1kMWBCz6PiWhif
9loxWVo1ATguDRBdAT5GS0pbaAXCMuo4jt+CBhIVNoRkUSYD+SqoUWITnLTfUDMLHSOFCm2Xl7BX
h34smhtU3VEzt3NBuPhUs7lLVUgWbg31Q5uhBsP0MqAj0+dfx+APZ8mT9mZfHu6W8E/4IhZdTHbR
HdsSwmaOihZRFpXy940VrdJcON/W/y22GmrMlJ2moSux2BsAYZvuhFoVsipoDMBoiMopUH3Cd9A3
e1eHzCUK9WTdsB8Gf7BK4H+5VLrOZ21fg8PggGKAULiT0gYTO6umLBJfI9xy8e2kC8t3tdZg7Vep
7WMVi0ZfLIU104pLAxVlO52Wox931k7ufPsL07wofe+eJCQQj5Gxe+ra6ylruCIDNCELTtClnB8e
hir45W3FHqAIwE6VwJNLxX2/sWCezIoFvwN56R5vfBtHOg+l38S5NOxJ4kobeAn2v/rHbCWDMtM3
mQYKisBN1D83LzhEOrAXbnENZyH8I2tE520+Yv0LnTOzdxElkYLRIGceVzE6dGZsgJykp+QM5LOY
mjZYj6uun7wZc3sYp3cR//2CvKPRPbWWnU0BIX1wxCeYXulcSVTBJQcyUCLombohkTzJGn4iHFv2
AnxG0nvc9mri/X6U2vyokGSq/Jg+ryc0s6QoVF4ryo09PH496Er57AukbTBfWIBPuMg4I5taF+3P
Y+Nxg1jnGrJn4AbXiw3i/C0K3q+i+7A3Habv5Uy1FfGIsu729jVBiDJbJ+NKuj/9171nSPDv3h8H
ZYSlwKlKWDK5lxSS7dOVnwzyY+bDwoUdn3Qk55P/nk9XKDD/4fHcCAAD8zJIlFws/3mNcawgvJ4V
stb+Fe04e5TF/6FMjk2LP9kLp27hyTz1w18/Q8ef2dooXdZ59HPhWjgJKFsnZC5uzlW5HCH76SGi
Vmx9zOexIHX/fk0dpeumeTzYHemCJajCi6l0KAE9p8wIBcNd7g9rQN2UAMsYfCDe1Y8uOm9L8xS/
y0UQGeiUZuvuuMJH3jVfZfb8wbTFJMbEN69+y/qvFgfOCDUWYdCnUI5IsAl1O58CJZxoM+ABmbfn
NmzIzTgTbUF0O7eQeSLXsikt/S0UYGrwbeJdIpUKgSmWvFTGTfibUdd1dXjknY2x0P2ZjFUWJblG
BcKkHT96tEccf8PwfQ2dmdjuXM6SFI8nQvkk9wh4EmRW5yty/McfyXkK3qTD1hRlgVsC2sCPGZBC
S2Dk4QfenxCrOqaLOO2+Ek08gRJPYSXUJ0bEE96bltkW+AHmf5GFiXdrOqUwI3C8KzPdwOpRIBD3
PZOj3DC3pO7OiXvxNHbU7zz0k2OltnR7QUmzWsMbaPjI4ud6MN2UC8MJV8pdXOwfzdk4QOs8kbx+
pnwLwv+0Q//1dMzwKBgpCF7CXk5ZJ4vxHORPGI09nQBnCllNuHsm2QYipPUT2pk+4FeyLyeud8A6
rxPef1yES8Bg/+QxkJPpI/HkvWIoqa36tHpCk1lvcLmgsrTeNgRmV6uVdvJoqsYeM3jvXHpCcWi4
CmHyJOyu45s8C9UDu+MpayASXnPYuNRt2KrrXY54Lf3OKemwAmPzoPcFsiug3KaIfomSZ+ces2fP
pxftz9RWumBtg6w4DV+aPJhnUQ0tfqFz5QK26FHERDo1q6FYz57zf5x7eg6ZC5ICj7omjdUCmJsg
Sva5uSqSuUeG/7vtDp8DyYo3rOl5gVkDD37E7JW8TP8gk8FSYB1EdA5avO57f5JVvYloHn3udaiP
W3pQrKjcD2rZe/0K4HAhZi8D1z7oj2hRIiAlh34NYu9j5Jy4lvUwbyWyrw3kbIwA1W1F/QmM8NMY
UFincXJV6isAlpu+LMYm/u+ae8Jn29O7SKV49I8G6GhYux93NpX0UZFzc2pXZJohasejg841WhCC
87hVG+TJnM39FGNOwJsAF7TlZislz3tqI8amF1s7JPCJNrr2XwzNTfg14cM8qn+fCPLD/Qs1IpF0
Rx+nYco5Cnkco+87XUl3vqQcnf9+fdxr86vVtrHtjGh4Uo6vsbOuBB6ms2iXqURtfZ68S4oaOU2h
FircW+QxtWGD2t9SkOtu2PjyyQtx1xDVsxd4sG1GGvxYyAhPYqhNEw69EW2Nha0dEhcPRUZqYPdM
FqLLbYbTo81NSYfGYns5CgEniBlA1ERZ6sG849uP2S/JToHzPhskoCx/T6xvvlkB5dmqfyInLJ1m
bHWrdtCH06rwqTudJhhu3qMFFOezAJA1uU7cqvwR7qO12vvePndRpqE52gh4qWFvxYLSy89uwePL
PTgLnpUCKBLdLan8iOhoX7MSdEs5gbsXhv0pCPykY3X4aWTTPcdP4+UfHZU/lSyb7qs2CSwvoIFL
Vy009aQVTdHq14uMKqsedx7NnSA8omMXVd95LytGR+w5t4y/IDxwF+kMGdDSZnObZeb+jS4LZyf8
434JAzR0HR0dGtnpDWQITM95FtO6rVO8d4mcmUXPEKOCVqvEaOBUa9Gc37hTzef3Q4lpw528rB/P
WYtWJP0uyuGg3RGyXfs655NOTM9fKcS3e6SKLaj4nv5NHHe6n/HrzsNxC43vi+uvItohOsXnFaho
jaN/xFJXTBfmoFzR2fTYUob+Fm9NVhqPnGzqEMh3+k7+MRa3PGm3D4AriLM4yBrpGaM=
`pragma protect end_protected
