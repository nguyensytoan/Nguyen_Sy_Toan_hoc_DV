// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:32:01 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
O/eagn2M6vzMJmA3/624aVZ9yzM95OI37qePJlRVgZzn/iWQuGaGsHTHa0YrtnFz
WrGTAr12u24FHLBlxHBJrIdHHjgCOfhrmnKGSzaz6XjN+aSQMEjsn4hLmew0r7u1
+50e8qWOTFfXLWtwJAZKjuf+quTdRVzik+S7xNezeQY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48944)
KekuTe4kX1PvnTEUPcU7ZgtNf8/xY8hJ+6zO+P5HSQiJNd9w2BhoKJu8oU2+pcf2
1kFmcoaONlFA2UGA+4gRsLtdheLZUIWPL+0WLnS3JijTdKC8mJS5D3M1KYiWU5tH
fP05bMs/kr2Pa6dZtxJ7PY6HcOM65S8gbL0S/7ToI87/sfWZVKMSr/h+eXUcW8n3
KfMr6Q/oOqrm5+kbrWEjjjEjY2tIZvjzC1NdG3z6OpU/bj8CZa478r9LqDZ/Tb0n
6XXJp3b3hr49QOsmq2X8CrfJ8HwtWeOmk5fpi7mjqBTGVw9n2Sjhvv5zJBg82uyM
pRjxXgFeoSegPAN27GePMli17LUnfwApnARTD+9EK12q+5teq1iBOc2ez685kYl/
7LbaOtdZPKef96xq9163Ie4fj+v9v4j2RqO+Ss6qGNnVBmpUMsgHQQLmO4eK4zQe
LvG5GhYE+HXxtOVD0CizL+VXCK4c+ndcXrNjJScM9CsSAu0Q2LotSN/Bg/oLu/td
MeAUMDWIQkQVjgUSX2Sn/W3i71p8FupEExuBAmL5vc5pHRjb7D1c4nAFIzyUVLUo
prWlf1XaZk/nTWeiyW/egYGdlMK2B1Qi14hIrM3cgAQiHG7pZ+c0MEhexebWLDZr
VMACdEcn0Mt+NPsnVV6Iu4ora2pnZAk/OBfRenrGABGCngpd9r90hBUECBW6T5Xy
tem84V0h1l1A2ejrgc4FjHC84LV0UkmGhukZtW4goDVXs4VaOjY4/KyKBJEvJmgT
XXIV0WRqW1JNumKYIDtfSPY0DFEavlgKdbHeLnOyFIV7vAN5nUIAJVKdzpDiv/cI
M9swuyWgIQWMdzY2pRP7cwfEu3oyAG91vCWNwOplOLN+nnnj5AMNenLdaPfvSLyE
0W4zx8JXTA3cXXe1tphLc/w/YEYRT+Sgql6Vnlupkc0QdbMbOgXhGpxuGrZFRTdL
VNFZ7sDyXaKr+wObovQQt/RyFGZgUtrDbuBpswWIMZ4huUfd1R9SPvyOkmRgGClj
1PoJ8Xr/z8eI1rEpsHPGeUNmCl/RZZW2kl2pqrF/eWEyqHQ0uTul0SvzvPHahQ/w
eHUhtCE/y4kSMRg1RMUqwozyqDQFhEARw/M1kPHEk6G1tlkGRzFf8rrM81wAf5ko
+KmYFWspWeXyLwrNGqixDta16areD9zmTzWVVfh0CgSqqNUQEmwZzmHQUYCe4cd9
KKRCnr6Rc0nGBiWCecrpJiNfvtCgzYsWvH1qwPfmB2eIosIc2VEzbmskKglVErwa
wd8LFdXy4M1SQvQ98Yd7KmkI90HPo6GlC0cnT04Se8FyyozJnILGjlDwF753aEvv
ATcf70W7FKWuBQ4Eg3Jbihfi4fs7yYhC1phibA+20L3Nn3XsfQH4JhtNI4Bo88E4
uhAvN5c4Jk6PomnMQLg2540vbKxu47+oVagGHAxRHeik4gH/Ad0wc5BXRYmwPgX1
AarOHIrhOvzxzY//knVF7Tf9MJfxCblZv1X/dfvreE1EdUPW8Sk3FM/gUhkmIwMc
So/afhhY5Xpnz8oKsrYhOhU2RdG0vEylEiUSmUfmDSNatdysT5XOjqJnk4QihKCB
dDohNdt6ayb6LKlVkRq9B0T+YTSKSZJWf4rm3EuN/gr6T93pu4I7FpQfC0x8mlxN
JPtP+2W66g2LSvXt7JjNVr+YB5+gmIjDabc0rd82cnbEctYxuqiWec8RXqXvICpa
sGHpPer92uhMsP5AOKVfOFHo6BEMJtC9z7G2WcnzmFLw/DMmGFxPpupvGQuzu2bN
+qg1RS2+iRl5PKHS9ntQzxFYrNEm5CIbMJ2HF7weyVVPhwIkQoLzjb6ReyG1GhpQ
S9H716uaZnFnGFtv+PNw1Micc7qzh1qqPWr+CmQLzsQbXlgt02RHNouyUTJxThQ1
XhKqz7Az3zp+INpnT/bmbQUVMRyJPjPZ4OafWOjE/CqYrLZkM117RAGIBXm2XnMH
Jj3i/XtVIJaT+WKHHTjtCzll6AL4J2O6CLghnoiT3wr1xAFUoF0w1C7TXRBP+/JJ
8uRNupWvLS1r5Dhqg+vxaWKGRo1ALf1+nNoQ1nMmc8Kf/+OM/aaxh2HBqbVwg8nx
JBGP7Z59V3McQT5uTgP36kqmWJxRs5ZLKpfawRuQpfD6KfchtZH5q0UD+VYLMVlY
EU2PmF7PHPy+gTPzmYF40pXZKYdpohx7A34fcEcqCytgV3w0yZraqx1Xzz/lply8
PP/0C0uj9sd7h7qqzwDU+ckq/4/tuuJSSzANS9rA0TPD4q/7DgvBEvqvjiBSSUhH
yuPVymU2KRmop+Bt5UmNn1Tj8hLtrZtRZMqqYImjWEz5IbTQbD5KeiDU2fIlD+4c
87xCvJ6q1/0Qf2+zn+HPtkZx3UA1XkklbFcxxldPB9SL1U9OotozleXYWAMPK2qT
JGj94u+mvp90zkqMpJZvoP0R3kdF7ir7tP8az/HbVzOenotQBPlLvM7yx5jqMTnv
ev7URwRC7YB5gkARgMKvITcOYGBOCPdYzrjejq8GPN/bcxsAKA2nbZkHbowxC9d5
FM0KwGhJkbmLbjMw6CAP12mTWx6mOtE+YUnjtGStAgVW8A2D/RSCYwUb98xnqB+q
rbCAB5/iYFgZvB5e3BBk0zWlh3iyI3/Y9nuOdDkQcFovGvKozQxQvRCSB437PrND
5RY72wFrtNF5G6+/e7ZiNzHDngmwC+FamVXcWZRz/dyYUke+0pHMggdkhqYZwiBI
unLZaVdNnXYFmu+bckuKUflCJmphXOWd/v7c9lC2edbaWdKdVXOtCP/u4xwIjeGn
MDaLTU8fqrXfF8h73/jRF87WgI4EkpvF7TI83+FP/lCYib7I60Z/W6mPlOTuHtTK
qVfXBCVT/XYIFcYlbWcw9L7Fy5Z7gYqHQ4cz4vE+QP6OgYwf7F32jp7VWRakhz36
rHGckmtATIgK2+tdezg/R0iJJ06WjsEIW5KPBFHZGir+2W/gy/QsIU33ODVpU8ih
83RZU+z/gKOByVJI1kACX0KPb6BO8xyXUSYpbFUcKx6UolJAjnal21+mqAc2rBrX
ufR9Q/J3740UXLc1P0C+QSHYMguhGRsLv6OCTtP2G6yAKuJpMrED5gsoNrlBRraM
XxIqgyvyaYV9IIfrf2uDECd7g/YvGLzaJDCoBYK9jqyfHvsFk2l1Qmp+lmFMQ38l
wJWHcNLzldbCB7eXD3LqEHm3ltoNKeKyg9q4PMSYC+qcTI9apOzsk0OhC/vMaubh
VMacGTVGA/K37c+o4i30QxgcUTbM6zs+tksx7ZnrmMTVNTe5mBx7vkcGafjFUIq9
RU/azWnadqrPimto0+JlfhNvYPHGitLdf7PBWD2IoTc8CMG6daJgSo/sMQ45D5Wu
rzE+t+Y/tP+dwIqtiaCC0RnqXAjlQAjGWdrV/AlPsOUpWr/m9osm+VK8hUkWzxB5
u/tmwAV1TG/NmSBsxI8uwqKN/cXuUe/H5CDcEOaWswaP9mzKtA0xkOEzzPRO9ky8
ltY0xin+NgApxBKzu7RqySS8SXxtHubG/hsFkW1lMeCUVAtdCFFtOAZTWbsjkckd
ohdyd0cts3QNSQU5GnZJMYX7qbIL5EENysGBRFf2cvMM2kxD+0HNdJny1FCY2Wxw
KnKhVlMqsWlqhwbEQJzS11EKyr5RgVuCMTBM5f1mUk3ihvbIKwDZWeJsvDWHOHRh
ltaVaEaAdgUhGdo8O1U8NhUt5bBCNtqveYbcbtmooSzTkE3NGQG3AVcAqMHazf9n
rqGKH9CGf7WYhxgyjP5Hhs+naXays6+LeAjpjeoeU2YEY16AHv+HIOHgle8kmRmV
+6pKR7Kx7u+llvyqWQzUaYawtawj+iYBLmuXN+dDEqR+WzADUnaK4+ICiXvcmPSU
56uld9+j4xuzvZUerF0r2fcRlvmuD12W3pCVoqvIhoxhTlhplSZLHSQQC5J9Bjn5
NMRKuZjZblggl9ZcOmYf9aOR3GxRJrIXyDFaT/5Wg81IvKUFJ/aoyqjbzRNpTr/b
8KFaRX1do2W5JMHmpckp5u95KDxiQ3sXH2hlpAC2pz4FcqYe6qTnz8vFXMGCxBS+
GehVqhUW8RedzklSg9AZFuxQYLDvm/Nzx4f2vhVvD3zOThx4yP07Mr3qZ4mO2rso
7icXYKTeKE9vf7vO8o1b8cs92dcxYB8R4PFHwEtN01JqdNiNOUG6+Qig/4v5FG+x
Z2VUGK46uYVUI99Sg2+/iRlmbsg++Ps2CoKHkqFFv56bb4fDgZq/8Yx7G/pJacwW
2/8DXuH8Q6sOXcMtSjt9UgWuX4GiRaSt2QDMmKiSzflMsrPIWXUjke41FYF4mDQs
hpVgSHp/UudK++BKFFY04D+GcbaEOReYaBw61ub72Zq9BD/UXM/vC9zZqH9liIR+
xw2mXSjUOv6xAgUJjqiD94mJ939O3w5vGBSdewlAk+NnhVB2v8FT62sOiTQAaHW+
OqvVWFiHXwA6Z0+UMhYZSq/q8FLGxx7J3rbXbvuhNlRi/I9YtuAYzyZEZ+CnkNyn
cCEInvkyMjtCoqJwtmbga7Iy9u3VkDdeuvNLTXPrDqxye0tUOMurGsf+C1DhjYWO
tomfnMtRip8ekBpQHUM1Z3u93ZioeFzD40a2m4R7SaEfPqpOi/YElghI2Gb/jC7s
B8AetL8w0mu2nk4Tpoxc1T8lDZ9JmWfrP+phXYspI4gwFNNVYmQifJf7AyFj1jMF
VmFuaUUYy2j07z/sHIOkbjIyv9Uloz1M1IrxtNHCKBhKsc9E6CgsL32FfiRgrwV0
6RRU7zKYNJifn8HBFA0wkEmRkiRelhjNYcI6X6pWn7Zc4CSvkYFj4ShejSVlAG3H
02OSZuSoXxYYu2gnp4Kb1E+cOny9QiPyYD0AZJFSkglTCvgoG2Gh5ewGliaWwZgt
0SD5vtlOb8SlAwk9NB4cXSyUN8+dj3gFyd3OroB34iorkZ8yWFLrOMbSsYOZSVj/
6mSvm1KScHImsi8nBD25z10te8UV0O+E6sQ5MBtPau08FWqcMgWxBuoae7CbOhk1
BbfTOa9qdTNFugaUjUPxxaX2ac12aXXdbXF436Yar3LIz/KAZGL/G6evbGa3SVD0
3t4WTmEUEU9MnxmlD8L5bAYE12zkWI+DPbaRNMIQDHGkHet/Z0muCgGcNbPvLsav
rAYhN7zntlExIhxviBamQC3otgGARqD2Ws+IUcdhRTITVEB+GVi6zOT2mBqn0d4w
lyXAIoYI5t1Od+JchuBXJHoRfXTOqjyi5L8n101Nt2QEhhAuN6vKOcFCl3z0gazG
2Iq8rZq8VeoWCL6RX/RinDHozgPnJie9u3DDt99jNsDqiafC1z9lbV5OO6sfOsEl
nZ/dFrfh1NJ50jBrcSRN4hngJ9vg3CM8PrkWdAt//2rC8HXm7r50V13QPIG4cibM
SaLnpvSdwzW4YkvIt8FHLe6bJfoN1yKC+cdCBClH8QdELITT9e5GYtalesrz/iMs
AoX3XwqtuSyFoYC6NK5+OvFzE+YVJi6w648GqocmUtCm0DcTmzQEbuwBu6dZp/0C
up54WRJ2pJcQoO+jGW0EoxFT4yi7LeDDv6X8rHV/Gas1OTJla6ldBCP05VDTdNHK
7VRjLy78hcWNKlM2TM5rLJre9d/uVwrNNHw2ZGVPuo31JD3AHlKN1/D9p0cLXMTl
ayVcnj247JahKhQ/8e9vZNp5VbF/IqD2OUCnls4Oo16Vtmefi62gg3MPpPkgIMoT
Uvx7ru7J3JNEiFLm/uIEFtU2tZVVC5DV4uPZF8AdGARkLk5M3SJUmF1jQ0HqnT8G
RgThLBnfLiioJfBY1WCyyLDLcIgLXODUYd4xGlb7DK0AobuB9CuiJyfboA25Kl3I
9P/1QydbCCvXYmRWVkUeju1xZxmi/5TELxBBxOGB0N1PrJpdfQQov6jCPuS63klo
3nq2IGS0YYU+CfY847/RgNe5aN+N8gmLfQrt8mIVsigyjUc8Eg0BtDZbFLZfGG0n
9OPW3TjkuahJ+LZ3t+N4vQI5VNEdgT0oZideu6mBSudmlOJLsqM3s0w7h0FJYwLD
D9pvyTB5npB2YyNbUfh/CUvCF13sGAkEY5Wcay17AZ8l4XA6foUD6gwJS4AIznhL
zS3vpRJqPzVfDhurOqLez55Z/SZxbj7ysln0yutHOLyMJBtKVaHQLy9FiBPcgR0G
Rezz2Mliuxh2CWTGX1E11TRtIf9dzhRz5AEPYj9CaD7PrEDpn5VMLIv/+RoV8Shl
m+5qW7yiS/HhRclYqsxFvYxz3eGzkySlhM6YDJRDGbzGwnvscdXtr11a3vGom4zI
H4/zZTynnGJzkYppOn6esnyomFIi3QCM0/jLiCgujmcMnhs7DWtGyG0Q384Crqd2
eh2kZrmorQnQD/6Mkgfu9qQa4Upte8NLUxriLK1Cf8DrOyrL+CDxyVnEzlc66ZyN
HVh4Y0YN+YC2jTOuv2DibUPqbmxSziZMBP+EkKYyOWUnd856zqHkyRseQ0puawmq
TiJKKq/N1SPggHe1Oy6LoAs+nhasMaJdsKualOmwKOgOKMxIfeuP2qwJd72O90Rr
9osEhtFB396UQM87xqQBWP3K5vGgERL93ugT0pzoU7msdvi3p6rO/1KYBTfCO/i2
nOuC6Ahft2hO6GYynyWDv5B6V+visvNHoh41cyEDzpqf9nw2rZeMxjdnN50wV6Zo
SoOKyuKaXEnwZvlQQANXJ2dgQw+oUMEr3hIpNU4kdr4MDGTr7alUeoQzLf8r7E/V
6+iwxmWPb5+/i/L8XzHrSkaD/FHnDQc2YeRvocrRkrNp2hkWny5FvgD34PwE3wjU
xl9S3M2i/LTlHuruRybSCKXT8O98fXrtEAAGVEYqiPUJZ/Hgn/MwFMSKToqvXwKh
7Mp2VZ9hAW0MBrcMLNQrzYYPtihw8PYitmZ2JBFJWN+RT57xOte/xyR0CgNfzEVQ
T4A6pxZrqo4exYXFVqCIGKWtqUjJVkl0kIGvDrrqpmGzUItsoXy2g5OrgEQnTAqs
plOcCUkgj3+N3EUtep+F6ALQYn27T5yzlIW2VYZD/OsX8WG6Ge1xDapOacsLOxxG
2iByURkOMLtTiqzYVf7j3gcXyJlPlVjdgsYCf/jb1xZxe/mJfpJUKaYjkTb03Di/
8N1g+6ttjd/7YqDzANGTrix1pAKqaHyOIlorZKGOXC4aTc5gNMcrIg/HzQNv1ZKH
b4Vh9EZbqqwmA0rn34EgHEbxZfwSddWNck6pj4D1uC6azAMM3qUInsEqO74IAoVS
+I1w8MuD5O/JDSpaPPw/JiXjb2av6xMzjheHrQfYWsXZqbWjFES2xxTLiykA0ZsO
CNbx983I8eexOoeso3Ve7Q2qd4Xrx4BXKCiV6kAt4wlyQG8XmnB/antUZt5J+mdt
8GD3tjFY1SzWR42FA8/k4WGXd81neob8SSd/uDII9KKfPeNQRFRxTFMSlmv0lTZS
STKWIvmD4ra5V5wr6GUBQq538ZvaO65z0bnHBwhg4768o0laH0fPZOMjcrOdDKqM
nOSukvpnf95edfox81FWo8ojNm8VC1JvBB6AyHFNQHa7+rWg0AwFOiamjIIgq192
HGpLm9WcrorECscG5gqsRN4hos2Cczpco75oJiBbQRlTMdPzHMxWkI0GfpjX8lCG
xnwa3bxrs20qhprCbBCdLEpDYforbnoWL3z/eKNsy0fe8j8w+9vRK7nQMnAta4SP
sILU18PeB8tU2MmT7ObXNLkhH/bgYFLEZiXDkG3FmNg1JM6Qz+SrXqG/N/HfM5MT
B4OVLe5lAz1IY4dexnGBU6VpobXyMdfm/fvFT9kJNRwEtZAxOWB47tTa2uwuw/Qo
A2AXfHBcQYXqz45hZVOVOsZDEy+amGX/ke2iHeY/N9avKX396dPBcBMxX8SygX/z
Fv0KX8MWDcWb80ExZIxLcAMCoY/zO3jO0nOq57gZdVkxi2d+L9P9J4HvnokaIbeH
tk2VVhzYmE91hSJ8iZbTLOjeKzTJslmi1PKtrOMAUG/W5YWFG/i1t8A8DZKYwE/S
OR2aylRw4ueY63b02IGNO3/AHigCn4TBnn1EfqADuhUOCQG4L8R7Gq7DkVX0/Bjr
IOISdd4diSM0FtH9DhUeKwmnoo23nMhCdjamVyt8H9JR396b8oX+KhZRb90UaO75
xPTTpxjRkE9TWpk6YTZ5ZRCKf85Pl0HcN1C9XV514NwEkkXpwvPicQQSO83kQ4On
Zutva+zuQ/UOYdlVR0OmyS6Lj5DZtuKDMMpX1Gz1HEgzFq5ct1JUCOAGmB1SXNMW
YFtXV0yIGWRwzu6IFcoxCGxm/1ZE0gBB2XP1/Aih+E64T3cNQ4o1hV18m8PkIWeL
QaWH1pClUZ6QKR2Ui+ycfzTFhDW23oWhwSkAFXJ9Nh5Yii9wEK93V6ryHydmWAzs
lhQYTLedLu8urY7+wIPJnwCeguCxUvtLQEgUbe2+/CnZ8XRRKwtMN5dj5nt5yNF6
dGyXW6E9Xi4lzCs4behGkFwlk1zv7xf3kJxxY1Czky66vhD78PP6cj/wIMo6DkNz
HKxo0w2qfOA2bYehldv4ZBePAWnLujtYvuCla5q8LzTeB3OBN8bc1dpHktTgPN1O
ApNlDIbgvJUKxBtUSB5JaFZK3zsMMNNwIqA5vfSwTGwEQrnZ/S0RbbUtrBjOIfN1
HICzwByto+DGlXNclrOMdt8crpKtggdzTyw2NmTuqPmFW84uAnQ8wMyqcKgOAIT0
Ko0FXXVNiCrc6Z+wfpKeDS3a76OEA/gEpb+nYfuYo2QROZju3ODsE2mbC/zuGX3o
ELhf1rmwPfzTet6fiiXR9QDaywVcJlMxqETztYr5LKHus6QfxjeqH+ZQw4KwhiK3
9CRSL7Z8yJ3nqszbnHzOEyMLk6LA1tKSabpUr4pyvGRDPln9CHj0OEqJo+OPkkET
3i9w3C0WpRI8Iqz/DQEG1XRl7WnXjWEY9yNPC3nfr3BBiz1jSWlVkNHdLIrZ2Mxq
oaZJ6t1+FkTcblZTJsbBOrtXk6pvG9kCCdL6KXjWGuTC0fUibHzFiPl2Yj9ttfQB
hqx7MwMyT7xktsFrpk+t2gGcbBk5A8B434roa4+/H4LmpL8QfVCPUyC18D9Tm/bJ
ClekN1uLdoseY8qs/E3aPzNeSQdtI6+92IxumN5tEnvj7I8Shnv1uB2FrrMxOTTo
RcsFRtCqkp7LoConYLKKV1nGDNLJ6V2t2XihC+4m0Q/lrpc4dTcaDm7mjaPJFAta
FpPdmHxfKfZLhQopMfDZGgi728G67/B9XKpEAQlqgWI4PAfAacL4eAPy/AqB70UK
MXEXbUfAThbynl6Lo19LmXCj8cV2GbxXMRQPP7bO0dEA73r0gxiKUxg3lSWe3de9
zo07BApw0nDKW/ixSSL0LhaV/Llbzo+uEkMOlec2Iu9kctBCata5GYPtywFEClA2
KWp0km1j5vtbq1QLrSx/7jELEs96a9RTT2cIMgXh/sak1u6Lvf0KR4Bzx8bGftOX
nEX20chO0+F9oSaY3xzKnaGL1tWh+GoYYLgXm5MJdegmQ9oo4zS7y6k84tPavrRM
YcaAPw8i2HsT/g0073QT4ahTArMAizJtN1tn8Ak0CosNHME1Wj8HuEZJu2d4CEmF
vXGx3i0UEQK+4wul9zLiKM9kOjMefpKpwM8ytSg2ea/MgQUxjcJsEVJIDm6N3axF
f2p98ElfLaYlNQvTeIDaUufP70Jr6I1j4RKmwSjXx80CzuVIh0y9fgb4JrIsyXRB
1dBUyw2Km1+XgCdWzKuGwZ/3J9n7JuL63m7f8M748xgx0kagkA/14jS7bUNa2QSh
fjsV9V6hXgchp9eJajtWI1S+MVsYfGigLU8wFZ8S4t3LSGQ24dS2Wlf8qgfevPKE
XsEKfYeUnJxaLo8LOENgrT3kvIOqL4bwY2dZxLs2K03iGgAMlA6BVGDSm1cnjjSl
Y8UW2J/kOnjkyzNoTRZu3GTtrzanoGFDYjUYYr7XoohxxVp40Y6JtcZrvEKrW60B
wPK2ojnWER8rBPJMBXu1zNgaHPjm6Ayh3Gm7E0a54v4CSWKZJGDQ2Dl0CkP/SQci
NVY/5wMkCIVLOc00TWxQrnfGsBuZktcL/3aDa+1T5ZLCSrYso/mYE0P5YWJXbapu
1doAEzrCtYAtx0uXmXLXRLBSMEDi+7ivKvHuRlyxcEbI1SRbkbSC7Rl14X1dUsu5
0TO0F8+4lsSB5VkawxYXlLq5xkSeHBRkTdBAUz3EWT//yYufhtn7Iclgbj0Wo5vP
DCMe5iAV2F4X293H18CIqNWguy9rJNqrmPGKpq27NZfpZxF+cJyFtycSydVnh6Wh
NQPljp8+ycbBo1Ad6PgqpGO00wXjLEKvNsxKUIVaKyhTDGwuMCN/T/wm9bhLZ8Wp
RVw4pxaoSqvKn4P4aLTg9DiKQz0SKy+eqpQKYAeIuoZCNUkN8TCp543BbZDkx5py
wU2xeUw4qhy4fUrq09ryawpEEs1KE/xSDCX4U72INKKLUndmJaLwglOT+58KJI9I
d4wwAovezDVULldY/9zV/40TPq/JNxhbRqUPRic5ExRd0t6Pr/JDATlyVl2mwQYM
Tl+Vaj1YlypWeOE2eV2Yo+UhlUgp+SUEUsdEoz5m+yHnfyPK8cG1Q9YQo4+/kObt
2NcIO2WbGvnon84P9c0y5tKgMYcImi7xeAKOSXKShiGjUXn06MlWDOP8OLnD7g5n
uXpq9S+ron0brn2XuXEoRk7URVCUl6Js7Zfrc6GTLWZ9FJCsPGdf4wrNBxkMyhMu
vQdAWCsXH52yQhuB9ZS7aAS4qXuVFGekHdhD2J+A8w83NeQQxP3+btvP3paGNZBv
/ZrrMrClapLE3eOhClzBSwTAdwmfblEbLNKie4NuZ8yjjwSuUfbMFHCDjatymO/n
NhN2jLaoSysKisNYa6Cg5jLov2A/zJ4sHvegYYcnkbkijsXxMUF6CEgpj478N2O0
s3TQIiUHBR2V4Wz0HjwDrGJfxg23TjlbptGTVppglBmlssgXp0/Qv2+E7BLynggh
brdrrmLWHbVkdLqR9cmTdyFeLikBexZQg5zsR7AhQVHIwXDd4I/N/nyMOBtuzlGX
izIqLxFyC1iKBuCKX366zaR3JtHMbxoWyrBTTD1USjuE5/BP7LOnO5yzgnsnq3WS
RaF9WfhWUBwd3Z0YpFSgTQfRAdyyYXsF8QIl6mAboKWLwSLqZUTQs9uk0G9tRDlO
VAlL5dSs15kPT0C6UFKS4VOmOtHXA867z39yMdN1N15BpsyubaYqzUySHNGHJMEq
5HWzGD2HCJm7o6MQehxgf/t9PKx6FrZil5YKvxl9HO3aLITCkKPgSX2LLVBCBDnT
VpaH3TOLJ86tQovwQFNrhlEbwPdAhnIqxXcWkuKQpGb297mxao8llPb5f3UNoS2p
PF25nCvREv8CYn2c8LB3hVezNaIBi2KwUK/x8oFvodMysQ5tji2jewL77Oplf89I
LOBxn6xeWSnABgO8LZPzfEfC/rGBIcs+tDinfj90DJvWpdyAdbZZeXVuKeYYUE+A
hC1g1W1Mex2BMbfotZP9+/KabsgY5ZhLz8Emw4LGQPp3jSrJOprimfwf/IWSDCii
5WsHEG/CWSIRFf/TdbSAuqMIsZUTQ1hsfJpR3G7DUzaL4QdwShBA7laCJ0tzGfNM
/2G0bHkE6kEFQ36ezGxf0JZsGYGLdjt74A4JcrMvWBYn58qCd65nr2hzVWGFT3aJ
18dxdwW08kecbex4rmVdZq9DAmV5RjZpIVkltgo0AR8Vb4yCmDEEgmzv09nHbv5T
5UU2blyFDLYNPGAjjL34So+CxAsdmg2jGZXbPkh4czpi7fzHOijy0KGe/nOubmGf
MccWc86VbMPl2xTcq26VLxNTOaSDR0AKGEqOo6C30iQmbclCjwL6g7HD0eVKpON8
CyVFvdM/lcJSp1QqZR0JPgbERXj3SOOSGPS49BlLgcdfoYj8Jq0/G3emEm7L6CMB
Bg+QI4NivUGLBUsuq5vPvyMFjSFv3d8ZfCIvuqqzHr//7JG58xUGCQ8qmUM7EVji
AFaFgK7Tph79gWh5MKzB0ZQUUZlOchm62pMMmBmLVmK0pSSByoChASHgq78eV+Zj
Oqa8CirRVB3OLHUioAMAwHnCXsdAy1poA8jEwrugAclHE7JsqtVIqNuqHIurFVdr
+thVsoyWR0sw1mZ96RIrHftlkJaUSK1KsXM+3RXY2gIzHEh6x6c5XW/lSOaqE1/j
8PhCDaD8WR2UpiB7Fzikz8MGdTAtjGUGn7afhtj/pLj96HjnKpW29b8f2ZppEk58
9lV8lbxsadF2D+5MswE/qaB6CSKHHu9kkNI3LGCvMk1zJir1p1KVuEVSH3+IFfPu
0mRl+dVckgGM+1rVBduwFpAT0Ikl1vKKj+lBpS3H2T8nGrQTfrnDvNeH0aqNA0BK
ZHXitvNUk3ymwqPwfCwQ0uuIrSx2J01WpIOT/sCZNscK3a46YRriWIiFIAWb92UX
YVd5/Xxiw5S6z7E/GPbLpn0okFiwRoxXidbVcszzps+btvzbiO8ID8689PkHt5C0
2KAby+9X2qCuht3vPQX/VvI3S2bzX+JXAndaum3EFDHEQbQxOsvBOmkRysyp5svF
7yeh2CXugVcVuP9U0G0K7tapwOumlsjzIcIwQpcsXNHFq5ZG1FdqWhP6sVKPMuAM
UOiUow77wBdJ3rGOyxSHKLY2ahndlUBB+vxO2UTkONeiRxE6sRhTlEvI/EsG0B3Q
+wjgHDEK3I2v5zRADR1MA7t2yMpffs18WpfKrdpmimPe0U11GQqh9w4tXrwj54Z5
cGNWCaIxFc0uVO9d+5vJL0yWwZaY2fNV5c8xDhU7cpRlfl1xdJKQ7nD56ZCB39z8
JGcR6OY+SjIqNQlLdYCOFm3sTvvexTZAEFWzhfRgI4+d4tO5RXALtRkA7rFOUHD5
m02kGGbEkcQvotb9vua7Ax1mFzHoEcAav3t9J/SX715tuOhIarRvmBl8/owBQtKU
l5/+428g9kquDvynPVK/j8geGPFjcfSEwUSpKDn0kK+RsAFfYqVM9XwzdkCko1xx
i8gcHVT4OgAWfTxb9Xul2Ig4eUCZTzN2kF2hf7Qokqcu/kOfXfwwjSzfrMQ6xx2n
LHEbkP85Mi4malizQE2slvdKaWtPbBmuLioNLsUfezpt4SSKLPkfxMLVHjweuIaC
qU1Ka4d5EKi1gCWb4lSVTSmARI1AcXQrAPnFvN28rlSL/FcY6cSXK5ZX6oyGujMA
pj3N/v7uapt2oNzUq1NdsmFOjYDd4qWrmAte+siVRh1rrrya40ZF/0gH/zDad2sR
zmj/TalxDoZAvl8dqB+krEBhz0i2X+Ssk9OhcZWgg/Zq2p23VchzvMNqDvL+SU9A
t5vtm0IqXaMr22xY7Z1+GlOi4mYNng0VAkK3t+Mduu18RZYNibEghchkQO68f24z
EQ27qJ8mTzA3mjBKmLTi18wblD3YI0fCOfYSRabSLT8LfUSSgCncwCx8DvqvYKeQ
L2vsOspy7/TmsCCohzjhrvBvA3a8N4vc9qhPg2im5r5k4QEGqjvjBgrW0aa8P0Mf
M1g7/jhyompFU+CJSMJ6M04Yh2OwDbdyhaE02ta4UmsHrPwyJ/ZFoUhSwvw41SdS
egJ7jOUgQsY5BCDQ5IkbhYz5BeQeyXlR4YjUPQ1nPKUHGWn3EyXyVn67a9bHrFy9
Xw1DbiDO7LJNQKauIShF9CFgKeX24NWvB29IBy/zBEDkQl743YFG8VaEwbYKaIsC
79tM+x54XKqqfO430IF7MTm3GE7ju1li9z6+1Bb1um0P920GLSn8akSNnNswLuvY
Dx9H6zLsT9HAFSXcIGKJICTG4/e/vB4RY9ktqFtamZQg5aK0wUGnL3JSawNSyoN3
AgL2tcSpGyGB/tapZu08w/3goB68yaAPkmEW6/1yT+ksA9+0o7hWbdpDidioeRI6
ifmQXXTuCHOfqWrlAAEIEjn01e5YzefwIhLlzGy2JrizizrGjkQ6D2VjEtGfoBg2
CYOhw/z+kznjE7VC0YpO+EArtXdfXWGEUd9zwGNtEWIO7bSH4HYbdBZOkE9tWent
eYFPhOX+k+nNvW7kNRWT375Bb8f5xbttEcORsHNzDW9p6cMlVz5ZHHeexwIGwU1U
w9WfLVilOEe/PB9if1OHQT/iA3UWcOcwxXwA1/HlY7TK9Sl4jRjsoFvPGL/uvvRd
tDaFIHIu7IW8HjpcRFV2lQL8iNhU/3dsudq62o2P0bXMMcHvL0migprOC+A+Z9Xx
w+2kJvcZjclHj29ckhRmKZN1BEMTWjWNcT61CXduLiRYUG/QbucuuJcY+ZBlZadZ
tbXKItzENqPPqCuuCY2m4xPaEuZhozpoTBhFp9D7nW897faKEBiw9eiGPPdj3uNQ
d4joZIcHAljJKCFw0Xzh+MEduybhQMQfAi6FEYvYY6TX3mfdL/ies10wgloj/oba
dLjY3TomojnW1YPdP6rKrbq0BmTaYF8wxbIvnbyrJTN/vAH5cqjp0igZHmcg1dNM
XFQ1MHLzI7Oa0pV8OrZzlT6cu3DXeaZ93oxBlNYjCqcBTZ9rYpxfYi+UoX+3zAk5
Ww7r7EhbnlX+yngdtesIGjTvwBVhUGwDGqkAk8Bj2fZrUDl3XBR3v7Gc3yg035Bk
Ed82PpwN3Qw4Z1EzAj0c7ad1g/naZILLauiNqkCxLHDQrJB6d+LhhM3Oe+M5zr72
i5VicKzoQZEE8yW0m4l4yFfx2v3Qkfssp/Mzj1tsJ2b1eR5xbyU/WjEvMRtuqCzM
ZhIJbyn/4Wb70c/ZukaUzxk6WVG2RrGufzIyzYiPBoehHlV3UVLbRlDCc/OkK9Yd
4+S8NGHmTHKU3Wvt0Y7lLUVuMP/KMA1yt3qiyDZAsMicldhmk4O0BpALhOBv/3uV
9wHuNsEoe6XBgLmtwRrS9fLZ8bq89QYf2qKtsi+BmRmITYFVH8f+8Kjr5P3eKsMk
nBL/zKRtHoz+Gd2XtSFxoo0QVOXMkmVDx/wFQjB9DTf4RCOrUIOa4HGiqXJqVOI1
9XGVKmNhT1NOn0jlxlXw25L9qhZsgp0YlZICUz+CDltFtT704Z8HCE1k/abGTUgO
HMcYKS9VPaxjdBseGyRb3jIltNf4Em0wlE8/uPpE71j9sXNE3YllKZNeRIH/vpTO
JhO3sV3PWZGM43ULWflFTShvcJvvseVhu4ra3HpHbDkpcQhbIoerhKl241fy43UY
EC3fT1SYRbxEB/ZnGt2+wBNL1glxg02qjnheuaHeegvUpnycowIEG6z2tk6+DLzj
6f+CRi+475wDdX2qlTq5xURvjaSzWYHVhc6v3JJpKv88TRv/Oh3M+KbhmjxOp8wZ
lNIAXiq1Sr4ly4dzq2ZgjNHsLWYQAqEz/n8fo4yjVE2+dS9rEP276Jbvv//pIDSk
QD6wSZ1bPMyf2vvj1e6CLO8yvrMvGTG3qJm4Uo69NEXb1y1/3qPEm7qawWf5zBqD
NJUHZk7UrYt8+YhX+0kA5YD+p25ilXFOsE97ymES8foiX4fHQ23MDAoLR9zJX99g
C0seGCpXY3sQN082b49V2XixSdcypP9XHBuVhgt/8qokuMU25RLKgRiu8ZpQz5MH
nW8cBxOac3OKgZzB591cC1r5C4jPQVG/fG2A1DWapCuCh9VOTHBrLURwt8e1jdYJ
TbKpO1HEWPlshSIvOHONklq1dRdc8fm1AcZh7SRQAR5Fnbg8Z3S+3SM3z79T6+Wi
l8gbK7P8QOgizpOsKxpzNzgRJvK1jaE9ACOSZ0rEHAiLbQvsTAMEC4sg6shtA/3x
VJEyHgQWYWl41QP9AONvgex98e/sHQ2jxaYgEMwgRgTxpgQYww78kFTLVGNHc/9v
WQ+P4NkAFIBio7WTH9gU9E7P6iZ4cASagexNL22VF/+eAHLpIVZHMozQxx7tYvoH
h+oJ9mHUBJKsonQtffnSSHFcyz9xpvDQvdva1/dt23h3bbJeC700VdVc1Ny6RcDK
WmIrrsMv3XpnMVdyV9pLtskP/vrxNLKOwKX2HsoVYJuUpzA1fyiz9t0SOJtowACP
EL31phmiHhIQe7pwN0t7XexzE3LKck22fVOKmoEIr9wadaQ364mSLHdB/GF9xS85
lP8CYPiLNvDIwMaE0Smdu5/cA/vRboK2QQJcfX3p9QXTFag7J9Hvb3BEX4YEpGSe
Fp0xyQQvUsU2a4lU/bjLXTMGqC4ycO7viwYGj6+SKTrUcd040uxfmVazCTk2uVwf
EK9pcMYLgr1JKfNwGZTHgwaVdmwRyq2soTy7DqY637u2HJfGud6+9gOclBK0cVYR
1Ms5Co5Ni5Q8CCO3aWm6oMc7nOqrJGw2T6YSx+d8taCHqShX4OnwEkMJ1jJ/evCu
QWvuBImj0k7tjf8v2g3zf4uQXAiHiASzHNTl9AzmI5e9iXQ1CNRacjOKskLsFWz6
EaJySAZAqfkUGwBDDTl4YO1vjHLqn7cOFS1M20MwfLAmUj2HNGcEems3V9sCPUHt
KDlSEY8hwmMM0pBV56M4Dz8mettyK9DgTZ1wjCGGSY3qmwJqIqTYANpMFYf1YwF7
k53QP+360UjRJg+LMcYGB2bibomF4AW7M7YRGLRbMYI1ato7mlMduq3mstKQRk+e
ZQErNhOJ0srMKHz0bT84zCgRPkjqNQudOhj1zcFY6/Y0vg/deDST7wt0HnWADa6X
W6MSa1R0sCgaNzPOyB6CRWjld2rI6a8Y26asSx+Oexlxqem4BOr1ZKu/O3n6ZrvL
5EIVHy90rJdCpShTVVyOKHYysZ0tFOPRPasVA5TKySrjIxB6t1ZDAICQNpZony+a
Ib8lW5WagBkksMD7cksowiDVp2cehh9f1oPMPOUeyDI+zynH2eVa6RjgUf8PQh3M
icEysrRHBj6thOQFZ0hzHir2vMo3LoGuAbcMtWDwTIIlZzZTVZZmdPLq7WRXf+cF
dvI+mR7PbEiYltb3usHZRwZN/csNYLqyiwWlDIQpT0pE35UN4m0fxVtIvCWLrr+j
dFzxrZlBUacoWharTm22UBdotNTD+cKQboJf71HYaKy57R9opXfMbEy+uXg2OM4Z
VtTeFI7cl5/qm0m9iEMD6LBSlilW/6mi5CwEzqrDpOuvZg0woaLXHhDudHQtn8Cm
itbgKuoOae9VcJfTXi5T2qdwSl7aY/m/kd/RzwWjFy6PpvEwr138kGr+gO8ccrit
18gZTxbJ68gleKLT7oSIWVY39/FIPinUBaHhP0kUH8SFh2CKN9EdyxBAMYl7h9yW
CUrIHXOjYsf4JxU+eJpm1l07jPdFCrFj+UnlKNdI2HQWzx3BKHvAGDQd5LXnJS2M
3EFy6or3SkKeaqDvGZRZ2ZUbfmH74RUN0j31foIGdnMmQbc3kQHjAfstCPrRQJlq
i8toZpHin+J7oDqSzDjcaGDRYt5mdjQclJqeI0s5AVLNVJEyum8CTyYBa78dHM+k
JVlMyXviz1wzc+qMLEoR40Tm0B0UzWUp9TPOfemMYeQ66IyiTi5UPghNzNJyXYMk
1YqzvbgSdzvmWpfIrpWEei/XUg7JBJEfEOwurVrz+hKxv3pq+uDC2pIePL2Xn4Aq
A2gzUuaFvDDanA0FgM/7SX57OvO8Rh3Xf/s9VZf+6+R3JYlTglz81+W9Ztk9JDgp
hIOyCPreYXfY10miOFI2rFfxCTBuABtzOXW5PaOi8wZI/s6ER8BL2PB9k71Kqm6o
PX6gHFQbS3srXmmEopx1HzaKMNZpBA0RsECJTPn+eiBrZQOn2RxIpS44w8p5ejl6
+/2bw8YQcGzCh5PnwqrS280qF3xaIG9/MfHuP+lYM+DkPObjN5FN0d7WBFDuerKW
WVawJ4ILSo4o9dmGR+KuCMeCRVSSVxKEhUDhueBReEPRn/2Big4ZnDmHZBHuvbHN
qgzcAgnnjrpyLzqflTGsVDeugJ2T6FZKXk7MpssaQ+nDNE+RkqyJOEdByGsyF/+T
3UIrr+088G7N5xBxnFkXCd2Nfo3+cfIecp231S9gVifeyH+yaiHSfbwHh+MEk8Iv
Ns2hQR0SjtciGzEDhYt95267WB9lYlEPVmP6SLcM4XwJ7AIss4zq7pzaSq062apE
m7okiD35+9Ub/qWCgCOr5YwSx/ooiViyElKYD4BDmlxoF/ZGBBv5X506qxGo4BoV
u2fMYpYPPlkkWgwjami9rdXgS3Um3Phu5nF2oOoThW+Cr9RmFSx9JV2JSiYk3paJ
gQ4+PqOGG+fLYJwXScWJSN9TIuMNjQPaV56MBOY1rgdbDk43y713k8vRQm8qdWb+
LQytYr3WaEEzbfli8SthsKdjy/KuyCtphaj5wOUn/MQQgkrxlC+3mwRdaRRVbDQ+
cBbW2Byn+fBMrGZohoiXyJLpUUZAyFseJ72kcXBXICTc2f23hKuUYeJFJzGsF0lK
nzjEiXyIg8CG6QuJJUdiOuZXzqbixwBYjW4jxev9KgKTRSnDZfJNowFVrSyD5dKy
dBcg9VKNazoyacsxNib8qxyyfsu1cC5AGjvrs2WdJluZjepTwVMHk/TZ8AQrYZ7Y
bB09EI8p3xsbmBfIttlsw90S/JmIgGHr5MLaxZZZJZCnUhN42SN1P6MjGMOEQRHL
H3h7VZbiUavJLUD93/V9Dryj59ifq35cicpZnmx9z8BSWlpneakk3MPkQDEgAySL
nAmroFWYEoMVLh4z+ebCTlsbpx5JAPkbHulrkfR2820QY9TzDXC4mgQBhzeVJjNs
6yAtoaQTrtq6AeH6eVgJtBhhnAMgwh99jdirOizXa2rK8mikEQwx7wzq3kv3c0vm
Ib3anugFXKHBHb1KyEw9WJHlPptghgOuW7juc8HOLOB/6pKGLyLbq3ZtDg4Y5NNZ
o7dnfKimkTQcVu5JkTPAZirSQZLRZhvqi+JD1DW12/duOYGrMLj3AGbUN0oxBV7s
uyC9Nn5H8uPINiyYKLHId1TwAcGq3ArKFFkxkQzMmxYB/nrnaOjCkR7JlRKNr7J/
0aDtzyCU4Vb2wYvw///MNH1s9DBI13P2xoFw4/qa+7WAQpaunJJTbdSLks8wZ9at
fIDjT3mo7dlGhIsXBNXdDD6O1s4lYRs4+TPGICEsFGcGBvxptjdJrB6zVqLNnQMO
1Nyyf3WtiT16NL/u66E4TVsnTqe/syXLrZF5gNxOvxnAd8QYNy1QCfCLsFjeYlP/
08tCdRWs0GvtGD1mQUNKM0p2NLA7zlAS5+aRWsYTtV/d4fo2k52M+NUJj0ifxyT5
ksYYbm6dsmUyFr838rK+QYggHdYqKnBeVj/zv2PSsaWCvDTjouM7G3NFyz2ZgBlP
JLkz4t2S9l6/IlXKS5PeicNzYL5pBlIelpXTbCwsprBWmD7L45gl/HWuqBFuvQuy
3iAUNnXAiZMgMyw97qDj5hvRblVTKHP7CXI6P0dG5YBh8kP2FfaU7lWGi2mtEw9d
l7++zleMGhRlzB4a1Bw9jvleFqbAAfQKIbFDfwM9iz+liBDtEHbxRE0rRfB6bfps
iET9tiqq66o7zrkAJs4imrPfgUD248d9u4Uyz24e0KOAgfwwBmj0ju9n/Ct/vVFE
DBgjeHP7MIClP6MgPS6V3F88RzgFizQ+HuktWy6kFYkM3iik70Mxs5uUfBCMGSMG
E0Xob2LG+80HgFnnpkFZUnXsRrIiQMYxUnZ6JvKYV9vLSiNf45XkhjGx7ojOpBaM
Tpj21PeBjsWxqJTVyXphzwoyuO1cwpWr8B7IyrZseiVQmUkZUvL5hxoEn3SPV9hm
aU2KYNju6mURn6sGHGWlufAZKtrLQKSggMygywsuauc8pJo4BhVRhsy+0zVx6l75
/zZykJEKWG4NN4kZtjHWGdyPjZFBN0TDj8yupkz19tWHHzD9ORwPiKUvfJbZvPYM
7gD3LVz9sQ6p5DRhFcI9fhclj22A+ovt3j/334qAySpLBLle+0tkBFT9F6NmbDEZ
ak3zzUEkzrsl9Ub2x5avy2zugtNlyxRi9NzBSTrt2JF6YTIzLN7Hz4dqKJpe7ido
Tgft8K4zLnHlQ4I1ckVnV49IPMexDmHHe7TZPY53Y7dpLVm31RP/a/Uwzt0ryC2f
us3XypGc+ZE5nGTTBSnKwraQ6tckJPhjJqEzTotB5GkOmArsjf5X6+m7Wlfep2Z1
4TxlFZpy0UwDLoEDhLy8SF8oggOH0uP3+uXVth5m1Ft2RGABxqRCT7FxPwlEYMz3
mQngaulKajkCOW5J/O0ZlCzRYK/TfPzERcwRXEXuK+IQRR5XiEp+UcEnRP75biRR
5pQ7BH5Yb8MN3kWYDSPbfIcsgDJLDpizmk32Fyq3Tg1++RL4U6HOXuRuSbkjIVDU
dRnzWDUK0XsReam5HwY4pe1SUCWQKfIoi5MP2kYb4trydE7ebfIi5SYP5bzayqKU
z9xLw91taJI2TZGifUPdSpjQCTeaEDXJKsgD+KnYgJpBXQuo3tsAyM1YKnAKnRKl
Iav/d6h1Z/1T4pM84F9Cm6xBD+qXcXNcPZ7kVaLJVJHR5Nww5oO37HbGO5wNI15+
pXDCDbl66fksvL1paPuYugMVf5hMR7+E6Bw1nt6lmX7H7my3Fp3TA2wELTYRON4a
VFEK4OGKENZ8CWM48wh3Cx2L0v5B5EeNUDFbKDYBLVeaaLzNtx79E/JM5tYnF1av
Wpry9Rzor+EKM7zGKbQn4U/mERPzAiCOLyT+GGk0w5qnfhRq58Ur3WEeEbtj9qCp
PWb9Dk6VyJzLTBztv3aH+RJUTYl36byXv/XB4sDPJyti7tI9Dhfxeyc1AkdfSFFr
aF0dWi0td+b5R8WTTcVIj8tqlNegyhNiKz/EPycRmoL5nlKFazrX9NFbnPPZ8esI
JWTebuaBBhIk//gZqEBC5QYnxxBi5pWw/l3zuXpXnXxUxG65sUqImCu9Y7LrHBrU
L0RZT3gdZaN7eep+QN9JHJsmisV8seU1rDS/NzvucDq/FK/0EadaUuZ3PUtrHzSK
YUzljHCR7O/NVQteWZeYcesDCJkEVYFfimSXB7eX1vchnmchBW/eFkwBgaLqYpKn
6YAFkytK8/7SmlZLT6KKLYz8sXaI9bMTSr5cQzgSto/2v0eOPqFZRn3spNFDHOXz
AiM2fsmhb7SiSVNRBCDwUF+mdtKEeMaR5TFdNk3hc1AWRbFrtXOzUumHnQ1g2S0V
Y5lhUzqD6baWuC3HuuNWmuzgFHrmzwSDHuZWM6CYTGlrez6l4u98tFlf/rL9qVgt
fDJC1nR3NX+5VctxecC0PuqRqZ40szUiF6GxcfdgGN6kL1gKZTMtrjdpdrm47Pef
2Ilng+ijZJ1jgDvGv2HCCnJMzcab458OfKkHH0zcXwWnWtT46DS1WahAJQvUWdSU
/H49Ln3+U/0muuwN0ZzOdToPGfins8p2nbEJ2E5hIUS3QanEVim60XQIpRCJYX33
jx1hlRtO+xtcyVQJDT6gFBMijDXH7APAIk/e+yF9luYLuOhZpdHYbqeMxSHmASdU
zlk1txNmVjaDsfdsIldF6xXJdq371+j4vXwYMBECCzalhxr/xWRrtP0nO4TtEM4f
9NCw4BmspYMy2zKSspjIT7HswiXEW0KkQQDc3Acqy9mZCA7JAqEWXaevv64zbS6x
GuiNSHIWn2awhUTzY4UgHYXEkjB7okKkDR2GtYv0K7vVVfCCF2o/NfUw4BZAIane
HW/yfUb5LV2z7y22bPLtTyxvLhmg01r81Ww68Z1blosugWaR/Ds/BAQ9WBfCA2Nx
0L3tr+eHuOuY1eESYIspJGCw7ALWQnpnWnz27titMfrX3vRwl/TTkAPlPC9xg2QZ
EyuUEjHD+9ppDdgpfiT9pMYXLQ+3u7gBEaOnWdVaBiTpZen4qHIKC0g1kCTzIfXM
GacqprO7plmrmshfkvdNHwpjIQStbc1QosSdCiM4A2Pd+I0HSvIMzDB6R5Ha+pux
UosC1mRimvv4aP4JQkggy02LLRHzdMD+LDqhiyMtvhiQ2/6e7mmxGZpqor5m2pVT
rDUYOeZBPkIfAvJPaiL1PiGXOvTx0CO83vaIuvj20jLsNiwEyL95mFzN+h3HNDGh
qYCqWI53/FejnZxw4hyRx0aaR/GRhtYYCtkMjo0y8K53lnhbDOucnxEI2mTkZjQx
wk5GZexgSVRcw+xdEDcN7aF38OHafB57Wb+PMk2kVTdredrzPeV4ZBAZYM46Cquz
MDHFtXW/8TlmU1p4ej+IJcw3VdLq68fvQmj0A5Qpi6VjFfWSOxeJRuEXo05Sadc+
OTNBpcW/sgnVC5k+lAYST7HqZ1MDPxbIiedCWJMdv21wHpc5i6msw0ORxlwDw6Wu
xTAjHnvWp9Kduixbd33unLGGeL9qZvjEWW8jbpURVw2mrNp7bh8W9PyvuIwRmrRG
l9viAzo46pp11mrf8J5UJ7bDAhc0FUx/qQiXh37tR90wBrm0b1f23UKaa7IiJD8N
EGfATyDDaPvOIRaA1nH180uoMg1TYz1ZS3PRclzIefsNfIFe73UNWXtbOmqYIQyJ
AaVu40fiJmX0+OcA39lqZem+e/QH4s+QMB1UmrtQkjKABZCYEdJyez14hiV9+l7f
rkoUx0+95BqVodo7Dcba8YZ3vHqALl5Xs78inbNE0z+UrvU5jO0bI1ep0UAu7ISf
imC8NY+NKe4ey7+vv5642Rxju9UBH8A67jjPxh7SqZlVdTUsB2PNwdTL8Plo2AM2
My13D8zvUJ7CFfZeujtmeq/flgT/yeFa4nZGDvN71MZLlmwyCPDoDprwfETLfnLM
TL7Votv2FYupf2fhu5vRDGFlJaqGtymMyrknTdJ7qCm0NCKUAqS3LdnF3OR7RWMf
9GhY4hIrPLB5Raw0n0wnu57wqLrxm4r3B53rYQqJf4c3x+Z9K5Kvtf2UX1kEBBRC
ofFMFzw+7S+P+Z9pf3+CLggW3+M//TFjZuGkgq9N4Fa7B4Z6PKk/XtXwTPBTWI6A
whrKKlQ/J+A+DZMHvO+Htcy4aIZeFEnro41aey1a/cD4ThknGgrdgY2kvNyTgTac
NHfYOplNjplP9RAHuufDhYJTAezOJCkPyHMZ1M4lMrSAKRZb5JP4gjHlpCCCzTMb
kNHeb51ulna/AAtcxMemK+3rsZDdXcrxu9FkIg3xIM2I2ZtslSg+6XNo3Nis2Tma
6DRjoZF4Ln8eYer8fs5dcMvPoVYQdDyi1XtifBqrUwt+vsq6+65vpbbe390SoE7R
zxDwjVzWQgDwqvE9JxOjumiQO3321t1jperDciQlcvyNvEufe+6QlOQ/g/Emke6f
6CMakhMd/v8CHsEZ1CbybVmShNTpELewRs85GlU/IbWnRWNKuLWXDMU8ZgNLicOP
SPz3lZFO4pSQIFDjN6fC6EJiHZkmR7fSF0BhEpJUuDi9bQLSpaaFivHPGVzQ1sm9
8/MSTRBe3rWEzNo2ynBMJZJEWkKhw9XYlkF71erGuaRvnfnjfS9RDNKUN4w0Odkc
1svaw8KQIES9ThPY/G0TT/iOb4dpvL35qbtBvsHzuZxaxX+4k5C5p/wxU46OfSpC
viV2iSSbSD6pH1qjZLGEKZ1cW3/OQbteMpaNgCZZQ+eSYtCAgyX1FQ7Y6pC8gPRf
20/bsHdzvQ+FUxGpfbseeldnEG6lOtMD8dCU9wQkc8/Yt34pggfUBc9BWfgORCMR
IDfEmVglnVFp9CLLeXclSFmqwsfb078VSy5rCChMsmBCgTgNKiPltM/7bWwcwt5Q
oJfc4pq5FaA1qIqxIN4sJSfuRH2wrw/pEV25mpX4jl77bdtgpuYXJEjmDTB3WqPZ
CyJfDas/LbK53GTVwlM56Zc9rCDbDufblUyvdGtaccYmcO/JkXEBBFDmre0Tw4vn
gHGMjnw+l0+N65S8JwcEWdERnG4znWCUuSIlhHlhQ/Tpg1z4Anng5R/g3A1UHNqH
dWmjfH/rwH51jCMQYchdbY6FrpkubG6gGDjI13c+cK9frbZWVgK3yoaDHN4qdywj
NLS0RYEv+ZRgWBQjDu3NQpHl/UCIYZokS397yu3MsJoPc4xs9/XW7aEM2rvqkJk+
fzUY+gJezn11faSU4ZOCuHoXH+mJBRMxEyQxzeaYkg1S4/kRbuHJVfBN6PuAamI8
V6KRc1vGUZfAe2OBpKHxeZNIMo8XtzRy06O+DTyfHf7Xy1VlTjMPf9yR5tnvPDfH
OrCk6lZhs7FsiJtz2lCuSxyQTxd7K7KPMWMXZh+xB7a+y2t6p3UELBbAaYMu3DNt
8UfPUJnH0OtxR6EzaeWbeZt3iSAsq+U3hdoJsidoh5qwRIW4zeLaZ2J4rFCgCoNM
SF9cvFF1XqK4iR+4iDZcVlQuzFmn7LcTrBTUisnfmNoYc4FAf3mfIOXb9ksm18ln
+DOnyUmRpV2iScGwVkB/ih9Vfui/0ulPUcAh0ItkDhITYJxO5u6PXfpf+Xl86RxI
xEVKP/1LhXABGecO8JAbEgzPbApoQRkiVKrXW++T0XRP2Vm8hg4cn99hCz5DuTvh
LM37chdQCCBq5DbQ28siOlho6QwDtEAeQ1zO52kVLp1zccoe3CSUnaPDRpjWQ1sH
x5GQ7T/3A4uVNnyWllnxV36LEgrnx2Nw7k1TpJ1lBsXjbWp3DYGCoaedPMSPa0Fj
qMudECC0ia+8haAsRJkYdtT0IJUhf+TwXHU33Wquw+0BUIYLf3yRyAS6FUNbQGd8
mJCHM4PKnIxAikl0VTnGwQMBcnTdbo1i0/T2q5ff9dWYvq6Sfa0HJE+pSuZr6ZhE
IEpUVWOX46rli20MlaDVD7SDazJupHrYX87iM89Rs1vISEVNQoPNxZrlcH/04ddP
OmBsjAF67oOW1iaXqjbvTgDQmNNDMvnvBZB0Njh5jPEGb3r4Eca89z50gU5JOY09
F4mSw6MBOjpL3MrYfZkdbtHLGVAEwHWLY8lblRUhMc78+oDC17Bzkois2feg1/hB
eXOs8nSkjhED8dyk0Re/sRiU4RziKGm4KoiDaS17lTeL5RJgaqrKoVHAbw7YGXJm
xWPCpAJchvwXTvymV96Bzb33XdgsU7A97NyTcjQ4sqKBf2CNZn4Psuar0skam+an
J49j/YCcrpDyj2u+ArJSTYOFjsRlT9JIc0MGSh6q++XFo/veYnYakl85KWOlsKv/
inuZxTgWkATQoPRvCUBOzlBd91npMlwC2JONBs4z+FroCkh6hcIpZ/4N5Z0zJv2O
iaIV2NengWUhE7djq5AChNfvpqF1q9O7ST/WmqNvcz3UCShFsPtG097tb+x712MB
w6TXajFc7fTJEDVpxj5E0w1bKTwkpnJ07JuCp+9rOUnZf0CtDvXShvgfHDsZJHuL
pS9Vyoh3M4vJ7H/CHnXdp9U7jgsmFe3A1oiuWXefQhMSFaMsfN7P2+CruqeZA4aD
J8HysIQ9kalS+IyOqFL5YhlYLQis6KIOX+UwhtJz1Kj95U0ScG+aINzv798enCgQ
db6Sq/UxxxJA2G+oVA7BRYVXuz2SdY7YJfV5hW+6V6j8g2D+8YP2eZFSipAG6IJH
r/zgNPcdqUiFu0rHC9jLI4HQ+dJbioAP9rhcT4FAFf7leQShnqWMTNyFAXP7C9KK
QxhxHgPsAePa2PJIy37DGcoqpZ5I24oUaBwudCKMS8Qm8140CYeGlwbuvwBe/oyz
ool4Fo8/tzQsJjDiKMIYcpnnITL5hCHQ82N6pLzJzT7vqIzzgY27nTxp0LoStZ5Y
/G58Gnb7zGpcSw6q8eW8gRJ9PP3dx6O5YU61o7B23nILOPG1WHsxppJaJD2Fi+aD
CETVcj3j14QZ/btlTRKDbXl1FRfHGBO35nIiuDqtY7oNRL+/jwZoM8xmbNODAQUX
9FDzopLiYUnoqIhDaJcX+GBFO5QXJG7grizfiFnfR8bY+R5qoSZ8C8gkDGK921EB
U6P7W8uCQxOBihWulu0itcjD/PwoWk2yz4fND9cU+11GO/i2RkFdO4rWBPoXsaEm
FCgktRRI3i6qhd4nqMZ4HAeq/xYOCkdRHYfWSDTfB1Vzf2Z1G4UVH5EzxK65Ejw4
tdIANJ+yfWnXCW0ri6xCwC5gjfzhilqk58+/WzCwaNwGQePC2BACr5Zf/d+WGVxz
yGmX3Pl7jeqnJA6j0IpCT9BId/Eia8KxzNvWazsyLIR3S8XcAq6WYcy0ALHkh0Mv
qhAeCd9oPYk9w0c1NM/Xc0fsuHATI4AId3AagrsGMvHq4gurGcSclk1Xxy4LtJ6l
ODvmbp+87if8/8jjDtZmfCYvkeEIi9BvS3aehdguTWTACeGyXoQPPtzE8LIxLWIn
wkPKzuESpAv3lTnZgrPChX0D6ABoMh+Tf0MYb6xesESwtzkH1AAp5JC0/1/R6IEz
F5GGE2JsbNOtuzvz/6h2LoMnb6k6AKXwcAMh04Qa3zNh8HnfbrL2Hy8U5Pxu+ous
G4Qb96lpDe111dtxPE8Z9FK6SYmo8z7jlivjBnVAdR9aL9/vu906c/3AVfHOWE+i
6L+dqg/Fjp5RUY0QSpHbe/IYfJsrudl3OE8UIJS3TUP5Q1I7w4+oTKPTf1ZcIARe
S2WS1l/kXfQTnx6oSaxOvJANWGWou5RBIZN/qb9II7OZAh8RX8/UUyAu5h6UzfoG
8Q3K2iCnyEwX1NnYHW1QennrUJejxA9WCwJGCGv4E+AEPSgH7p5qXje0cjqEY1Ix
o/PXd1VG1Ihb8og1F+8b7nBH0nsEh/Dyr+5+twDMahwHcBPeZRUzasLdd1d/7y4M
51S078w2PppdwKQUyrR9bC36mRBksrs0p6eh6wmTq6QUvn8jrZvVao1GScGhc3AM
7uPZO6ZZRFa4y5zymK6qk5yWYLAp2czaoAkAnOhzFfiT6KYePIylu4HZ/H22mNZh
2MWpttNhoDt3SpykQNFASNYcgMYcKdNPgwoYpDaCYW+MDiB5heyp5SarulM/4fA4
Jl0HQq2e/3WDdjw4ypNI08GT0sVcjxIJe4n60c9envSOAjQezRjuTTAc/POoliV+
J8odxekl4CFMNoXAicKCQStSBq03BJ1IHWFSnVXxGi1VbZrqxEmFuYc6h0rvDtBd
w81+DUXp/H6GmUCcTB065CG3RDruSKcGgQR9glQhKX5u9XbU2wwAKASwPosgWdsZ
5oQ7UV7sz5mSivKuFiQGgXRW6BTN5jnT8pBXIvSfrhP946LF89yhhNEKlGJzFRKb
VujPMR8FPDQ29e9CX+k3kuU9uPim8xue92Pg628yLLn6QaAkP/rt0AyfGoxQO2+d
kOuaJn+StVQB8aUDQYdLTo+Jl6C2Ow7ebPUcVKcFzXXNskN//++7XsEGJU0vDiC2
DwZnYmbvHBZxhYawA47z+ZoXPlNECw+clSDMovs6MYAqMommdLUvllxHk/63Xt68
LMtgG3/sRPUx5dkKf6djKc+J9xMFivOKZjBoSoIrt2HrAcxiPbrf167B++o5vV4b
udDFkgFd9YxtHgRTsFOrWhFchs/IN1yELLMByhof5jglpgGQBk09/diYdPo2/LYL
vGJicBkBYzieBdp8Ab6Gw1Bnu0Inu2zEWyCX3bboULnGySeHPtQugjAdkBGSOXeo
u/JaYgn5sNs+OZTJGGlHwpzu9mxvIDMLh+bJeHPb6r0Q4SPVdaiBdQZc+dQ58rsd
KT/aY+quW63Knsja+nCGlL2WsIfcy3kgwlHbchAUzLkke11d931PPH8D14I64PRv
EAiwjyv82RaJQufic3rUnkip6p4Fv5kQTbu7ODfnooTPfPEYxsceRsvhvqsMzful
zMxZRaJWSzADgltQpOIfDoVY+v/sbUn1Cfp5sf6P8NT4b8hpVeucUdqomBP/ihj4
ZC/BkBTTrjMEF94E9QR2OqzGV2VbFO56jp4pBHYGNdtQLxXRBKmhO1MLIngLJ0Yy
EMFU/QGwuUQ3rdLNmWjajScPiEIgIvd1tZwqkSvzkG/Z+KpdiUi822Y6qzx5cuhU
zl48aEWVmb0Rzcvd+yAHzXXXN3nGuNRSTcEmeDX0pa3PTUFNJ+Nj6NPLuwmjdSPv
Gc3ZuyAWd2h2sSViz1ZkYxXdMVwS4gcO2xCQrnorU1qlQuZCXv7ugPsyxvwE6ZIl
46zx23gB537ZJS/ZgXVHgqXZ6Jngo6xGK8hSg7Qa5eCv+wZN5rg3d5aImH7WLfZy
Vfnc0WL0T8msd80DJ8/eRyj2udm1lKoe3T6owmnecGFNmcpobSPHEcK1hidTunUb
FFyncZm+kNWvYtvnkoCTWx2G2iJ4Ro397UbuRxw52+xlX4JvfnbtA0Ol+XQqea3v
s6lWjx4ZpNMD/m1lRVLx4RB9spU79ZLwiaEq9d+mREcIm8zFaPtBrIML10neYePS
nGGU3sQe3aeMLXT8/AA93+mxfditPtHaz1pVONnP8Avddk1Onc0W6EVe5JcBvai5
Eok0MZq5Y+U0lV+GbIRmfVaprW2cBD66oN/nFe9ZkEW8CbKMfYBO1IYNeu8VuNV9
03OpXUlrNjAt/puR69hZSRS53Ae2L0YlnNtAsX01YKhipxrhMkolBuND34IIVk7B
8Agnr0mZ29Bg0mt9T1RLwA5jiF9eCd8mor0N9V2KP14EO0dE5VteSzp+D9Qd9vIw
D3v7nVhpun78PoJpKC2BVQ/ISutWuwdz/viGLo0mqSgHCZ0BJvp0rH+N24/3T/df
NVtvo1anSENnD1RmQZlELoHEQuD0nnpZQr4jwF6ecUTdGdgfN7ndw8f6TJpSKYxP
PQGNspU6qL8vW9zAIb3b12ZqN04wJ3Gy3CqQmqDOmrBwGgMxfSFUu4kM+bvw9xOz
pwPiQ2mIRtBXrDyFz3vq+Z1L5fvGVdlDRSVulQc+5CYGC4XKBbZVD30eqrFDvp85
Kwg6F5NyM6VDk7SSZPhzVPv3NCaI2Ltu3ORfhLh28FkGRbRW7iKFXJmBGJuY04CY
SViI1jS4J6CqNiqRWiPA+cpB05UNFf4aQq9b+8/AaEAkBx6rQMdZLGR/gykCGS/o
W5e4YnYpZMyHZtFq8hPy17w7Z3X090cWaJkttNBi/RO5sBcDSBqNp/M9nLs1sXNp
S+gzwx1dbjymmTqiZ3xPEAgdkx+dn45oz0Zl3AciM/ppqeyW6JfcXL4JiwuqOpQC
0Yrr8XhmeYo+UAyvM+A9UAJv9WoRJCsoGGLgNJFDmdjSkZjVzm+aI0IJnB+ghZFr
okDKby9nT5tyRtSP56euyCoF66fRAVKlTr+vH3DmEum4afs1oIGvtbulmpJnhryM
+dqRDTY4hWIaZDwWk8O9XfSkdzEVVNfwj8CzJtAj3DTzhmePl+2rR/BPMTVgzPlc
PUJHUe68RVK+EJ9zMAmCMQss6OC1jT5b7EANjBc+Wj7i/UXU0ObhS4MMPOcPYeIX
NXi1UPcZYitaFr5Q8JGSXWAgYPOOBMPuwWQgRc20CZtYe4wJwtuK/DyM+A0BoG2R
5vH+x8A19S+dCp0+cq6mLiQr9RzW7BJdnDuJvO96SX5chw6/SM35UCmvwtFEQPkM
xtG5OrDpCe++M1pZlWl1FhEKzxw/NoAfp1XTKCiBJbeHgw+dOH8GSUZZCpM9R3jY
VJw8tPpyxfj5rf1frgv5C3/InATBqYmnGYgrd6FVd7KC91WpYx3LXuLJxnx/WTbt
CKEmzQx2hCm9pgNu3E4HyNE1nog/ih0Lx93xHdpqO1wWshEalNW0BMk5iM3pdq+k
78g/2+vG4BkUe6Q6tCSHTg4q8cEWb5QxWYBdzIDuUvuhMXdrKRLzPgTwPLaBHGBN
saprNaQ1+PTJWf11L6g4UWQ5I32+70Mc5eJ24VMLi3k4qzQYHGjc4BKj0kivEcVc
3uqDof/HGWjBfHZGv7aBqHs+zzthrcbeGdfTm3gDPPNlJ4O2NU5FjbGPXjCfe6+w
Tmnk1mN0loJ2LkGpPOBQdtxhGb7vKSMtrP05ss056Hd0zUWZxvxM3lUOa9Z9LkGU
q3c72uEtUXC+/vSGiCAknLuHjSryiVmWTWvKM4y35XaS6KRl+P7Fcc2Od84vd/lA
MXVLNkbf1u/Tu5nlVqkkfanIqLqD/jBjVTIRruNCp3Nk2YTRxbFMyayUN6BmlsIs
2RUi3+Q6wFqrffQzv77AbfAgR2AzwEjWgnLoN96aLBIPCtM8WdDrn7M5gYhqbHPU
fxPjA9fr0vgzg2pimm6zQv5ZJTa0LbOqw1Tapk2ELcwdG/bywIg/IIFURC3ifxCe
6zsDcjMmOvAjWAu7auNzBOUi+BKnmej4HJdhrjKu4gIz501Kh4T82ADk0u3jwLGU
52liY7zk+4StJLijyxCsyHqWmrg/Lx9bP1h4K6bksfnTf0YbNWfV40YxYQwWn7bT
2Z6vcZRjDoH/aCSiLLI2HmAlOaGD83UOzG8n7+K3jp4xmE7URugSBuSkNMascccs
9I3I9c7YgTsfSPgXvNnAzjidAX1t1UDINX52cVDnpArIDuxREMn3MRL/rrygZDhv
CxVK3GRhdZ2S2j8q3jq8PFtbQxz8nzPEviBGEBtFXJNJKH6ELnyxN2KtuivaeOHQ
FxiHynqT2Dw7HZ+jKSXyTDETLkKya+ukpDiUS+2BgDyQVJJWLObLtm4aTVRdN2p8
yvr9T1hDTMdxqjF+qmbcuI0EtWEMLk+/xn0sIsOb6VOMAKZcAgvScW4WqkAuuDjc
uontegvCfl+j7/JaYcTeQXCifRQk6pb4oR6h5baBUIQQj5hv5GRch0ve8Xy8CQRq
q32JlvuDNnrlNh1CgVopT5OBpEb8MG8xcv8V3U25adveT/FyXF9NJJWrNX+8Mm0H
+qzOB8umsJccaabN3OWRa22MWR7D4RQHaxcaDcpM3rhFhqGDZ0PKichhVCJO59bC
u8JBU1jU4wgycqkGCLDgCrpCUecUpESzNAekKiqKxyjNlRkYiDgzsvL7TlhYyB2x
fE4heCZrZ4BAiQJ5FOVmkGSMlr4lHBNSoSNnRrnlVKWIyz1hiR8APo8O9G8UjPNQ
GMUnzJ2H+SK06BCNgY9quITJHt5BWFnal8GpIqp78Tfd4CRRh9Cq4rVsK4DBy5Hk
WFw1+qmhxblk7F1mkrPnyNwl80W0gUCqS7tOX9yu6RiHRHwrTorSuyRn5BSqs5e/
l1feNsg+OA+G8ulzhY43ZzxuN2s5nQOf8OhiTbmDaKDiMV7AXEIYNBB0qaHk1bCn
5Ubh+vP8jgeegc745S1sYiVFzoqDBDNnt2UubWuNXbd/4pONN5EFJCztS6wBe2ZT
nA2Zzf0lj6pB1MvaQ2/CMea/VcZDShUmZ0BQTvJsjxMelDHwHJ+lLbdqRNzZlOs0
AaSqUKT+uOORo+1OuvZ0SuTLtD/u3sDo2EqL9xcDwQj4A0UlRnLlGJK3XxA7CvCo
s4gI2Ab9turLlpOjs5bJ9T61zAOpCuhrWSmRGhw+kS5H6TdCC9wOMqCpb7FjxD4Y
GpSPGK2Zu/oHij1PjOaVhJQ3quDY2W+uhOsZMoXpx+er1SRPlRZNdDuK2GGhZsbl
VmHgStPDW5+6v2qIp9vd6VSWHq0YFHjU0NUJyBfZ3chAWxZB9YSRzrdz3blyWrb/
IDh8vDdzUMR0Da7XtJbNGk+9ejRlDWUeEUJtfRkHx8j5QsHITf6Ck2ee9h9iGpix
p3UZf/TyfzG297c1RWpJNT+9Lu6uVbUUkUgpbnXIEJM3qEHpNCy5N5fIGGg1QZcF
n8h7ZQUjX+NYzfx2uIfJSXrvvsFpjUIoopxyWWBqjvnDhUvCumkHg83mqAT54g4e
FJY90gxC/P3g20PGMcBGfYQk+8WL9B1icNrIfCr3gdaCGUulbUbMsSQsi6GLC1un
DosTLKL/6gzZh8HSdsH3ZGb1PsLXQYn9qb8oRdByT9L/mr3OXTg5zhZRZYjYbCEo
rbsugKAAow81MZh7M9UfmxsHMwQ4FXEmvUdD5WKtWAI/IsFekfWgLqteRAllbM8f
CbjDYDxl/674BMPv64NUerPbhc28L+6SLIgPlvulnauT9G3qG8ExwvcTlLZEVnTr
mD1NKjBJl3qjcVN3xpiUD9cfhyxK1Wxd+fA/ClY1ffeNCz9vbogTSNSWiGhQyJYn
bfuz2ms55OtHlkGmIH6dQZpfcpitvgLrG5onLqPchygL6fR8Mt69nKSVGfUSI3mr
aQIa2aB+djpdIxdrbUdAyYUqHgbrDgW/oMkPJT1/i4aQ/gScRuzS9VzcKbHa33wE
8T5YlQJU2Sni+TEcPji9aAmvLanxonKR84K0xUiLIRMbIal7w3qN5NKot+hCAsLi
PFzwSHB9NITFfQAyeWLS6d6ObRL6GSHhnvLNLi/KsUUMYpmU/m12jGFlsT/bGroo
s0D7A3dgCrlvbQ6AHvG7Fqh5AFl5JlEhBjpOw0P/3pfDflpLwKUn2N6yEyL/C/kO
1xPqcRXUmqlDEQNJQwgAT7qPnIXHFMPKolxcHDKc/ZyLBn0dDx5CrjtDQXUx1h9D
h6RufcUM2OFzGKt/jUgIhRKQ+E0HwjRKW1slqx2OoJwuIMxFAl0U/wF79meABou7
G/xKa4+1N5sL+05nlorsNafvOCU0Q3g9yMgVeE8NbVrZi6ZchiIUrprU3NiyCFsS
i0HmmdCLMpoFCpZip1dA2utjCHEwhLgbMVaaEzmttLojfsbQs51YTibzGfiVogx3
dwBen3LVikZcFkiPX/Kho1TSB6qJDENEpkQ7Qkx7RRsagpRCvzVd+yTQ2zpHBdBp
WJ5H+bI0EDoY39fn892poArsZi5vQc6qyVt4K+gbJreHGUjtPmSA668CG7dQRetJ
aktJ+VuhVdAvNzeh8Q8+hn7/ZJdhk2zbbKfPplo15Xp2zfZqV+FezEWgYIZGRlVm
QIbnvJ9SgrpILxQ8XkIKVnUAYb3D8SW97dQ8fUbE+DD4Um00qt3aK9WHGCTdsHWW
B0ATm4+/GppaZiD/1yhrNnzPtRxvo/mtB6vBfaHPiI3fJkRdhiV22XroTsXgaFdQ
WSNXEWvoeuGDU0bTnSZ+VWUanWGN/cAPIoxhmKstJ85esWmp4I1fzFP3z4cyqTU4
61s7OM6rXUrqNePwNA21gYilyRRSn0txS1OlWlFo0dPLXkHw2kKilftS0aGxdyBY
kuwJUujSWrmcJz1hyt1bs649dpwoBFUON1BdHrK5g0+nLZ/loivZe6yQQONIox6H
UDRKvnVmm1zuaMKGvpKFyUXgawV4KGMFSzfMsMQK91rwVFvTcuJn1ccf6j2E0Z0U
Wi4WDVAz4vkxTKYjTWWDZeDo+XTqpviB1iYDxBNPcr4UmaCy0UmpQBHZ1wPQLKgI
rkjI8KQ3yC1rS0IbGntLRwCdFVofKESzloLAawNUu52/q3y9nPoQTy3NfbLEdpQi
NgWLSApBmuhmKRqSy10kKWjCGDgMIjDXzIVuDSDUIUSjwB7KF72T6E0gxMrZBBD2
NX7L+EZK0xfYj5/LZLzd74hGw53LvkL0Ykk4w2WyfW0mLMe72KQaAEcLx0mkscOM
90dlvIB2DNbJelNfmAeK0Rm8EJq1+goe0hG4CQ2OA9IRhM77qj5H2AisMYjAZRKL
sne/rtGqFcQVQFK5Mk96FwUfMOCdoOOgO8gANGG0f8bHhe33W9Mya1W3Yab8I6LK
KKyjDDHNl4n13weIzRoKVzmh0SyKXSN821B0DwfI0UNoiqZklkqds4wo03qoCEsq
356tjSdVj/9lHkjoaHpvTX2gYa21bL2pb1l0P9FPbR8FAelMjAVlJpW//CiMH4ma
Std9a+h2u5LlBMZJOgdBMSPjCnUjmKwRpLjhH4XezVN8wy2mnOcE7GQoiWxeOuQy
L49Vtewgf7xZ7ugGFroAPsokllRJQPaRfooeU7ABKPB5xOJmPrj3AsWMmaoUjweG
8Rlbl86f/hEe4fwuXzg5UOcjMcF0AU2I6Nx4fzBbk8NDNRM2aYE9cKJR5osiVQ/U
jMTy0FgZ78ynEJec8Evkm/NXpuyxXzTQ9UNrIb6RSqJFosu5XEUGkEY3K/dDjS47
6a0yf0gbDr954dSnyuASYYjx6TsSDmC9byHtphZmJ7aOz7DAEfFa/h1d7/NveKWQ
LwDbvRoHxq6gASRGXGRWcKOUc2ov9/s9w07j39YUR+oiOlAgsQ8Hd856oU5Hck9q
6GQ4BmfMf/nzb3FUNPoy7v2VX1n5LW1NIwUyGRjBLuwGUEi2vhYz9+xpjQKFfocZ
OtFn44YNkbpbfebjTth/sxbYk0elhhlyaHkX7BJ39vSOp2e7dRuQJPkZt+EsXTyO
PR4oA5M48pZik9mNUTlynV5EVSpOX2ij0HI51Ipi7UXtcilRtu8lcwt8/RbWK/8Q
UKkqFlOCI8f2QupycVL3tcgOMRTAo/jsLv6Pz7OK+nHUWU1j92M0sj7ZWMxVNSjM
KT/23/qmEJsELA3p1zmFIr2BR0/JXKQjvNSJoioC8QFLJRvd0wgFMXwlsv4Wvguh
eJJeyuht7B/SSvx76PWR0gsCDs/JmeItDM90vk67C1k+WFxYL9k4vAWQWZLZ3iGw
9IBEiIPY2ypYL5WVQ9akrDICdOlvD6yPxsHQNJ29YN5e+c5vnfhaRYGlXPrlHuUp
P83Jp+abErI/JOP/2cgoqRRGWxRz666fqSY3M3saqu0NcfkBC3koPbJDq8AADZIh
pNEufWuX/SuVkdKP+4apjEePhnlj0cabFA1HGOokiTsDlevpo3AMLl6icn7TVm+Z
am40E2uAFL2TKnXOjLPWkT/PF0+X+KYF+C2dT6zzJv2Eh+qnKc0f84QuMlWG2OIy
HUdO/A03NPIuOzyr4fY3LcHHWc1VqweGL1Ipnqxt8r5FkXNM0VoJTSaHB+tmVGHU
1+WTYKr13RZdQ4N4H+QA61ZUr9gMj6DWdIsdjWiUL2Mt7RbIo+wJXIqCaRCcAWJ8
oSW1DOgpk2EGgqYPrSUtSkyD+Cs9E1XykzG9lsQaoX+f1UDPoofZvfc+jKVqXKb1
kk4BehqdLuASaeEHdM+K5oRQqRBZPO6xpjld0GEr3PSPJy/rCAVdupwPnxTrXt1o
FselNmFTYzNqZP+x5BlhV8o5cHRgc77WyDRGTapXNxOX8WCPjk05Nx+zLch7J7O+
zSgwJ3WGAnvsbFGlAW64c0PH7Cw+di1/NjX4pF988oH2oluXtJ4RqvWVIj8L6W0m
zUHZIn5c99e4f6BYUXdefsX6Vba+l0ATyp6JMvAd/jeNCzgxlsOgrRnBl1gUEnPR
HNpFj090mmghZHAt6brkmObCq4M+cTsxZTImC6YyKWEV5SFaZXkL711dHOb7RxS9
3NkRFDgVhJ0KvBIF3IMAB6UfmKWVtfWZL1FrOTv4Kdm9YSQ0U6ZAiGEPOWGQ60OH
HoyL1RjpJ6eXND6XOXbJqQDt952hKC2JOs4BId30sMJesk9GHsosbDrD2Slp4zvc
4WuAfqioGdcnzWcGkyXTfhSUD/RrLc7JtiPEwFcQ+mEJE/J8medUkxJDXqN2pHYK
Ydg7JnNTXGCdrbgK9Rlz6c7DS4R6y+JYjdsD5eNyLek0iHFJQ6aaopH2S2+7wVZr
s8OFmDlQGlRcQSA2vyBKNNKpMifNHHWM8K7VMGT0Zt5opQmD4vKnTC6VTnmnScSb
w4m588oPyfSB9KXqO14WvCwJXBTrDvQ+QispWoGY78AlPKz0PWwHFd5hZwNxslPj
hksyncVMGPvY+jvySDyNvNGakX49FOVM9mcLXK+asGT+JG+BFr9xSohjZ5Xu8fBu
p/jep00pD9MO5FpZSwJZl2rOVqKfIKzAtoa052ZTk7iW0cYi80iCwJyFZ/rlhOGD
VfY9ZUP2TdeOclEL3pg5X2Qftf0bvJXcTarXJPm+759tz7K72wXt57/d++tzY7Gr
JGuAN01APgbJMqUiLRS6drMqWcnl94OxjzLXaIFe3pO4kMVASbyDFE3PsGtbS1dO
q9epUoPJ5iWPa3kR3Hs+NSDP5hJoy1t/NJbTCczrW7A5MOMA9HRDADY5cxyYftkz
sXG2vNEPaCffpjQBrCKcidxKourcfU8ceKm1G7fE/hTRnFnOzL1IiHo93ArO87hr
oi20OOfxEknWtOXl8SugjPQGlWuVq+tcl76Q/SCdcsghJCeILGp1wxz0yEjfKbP3
1acYL+mfOnLh898Qpxwd0chixW1Xulp7Y/IOPFIy13y4mclFlgM/DoTtF9qAtQoq
9D0RxrCVBXtBk2SWuDm+zMcICwLKaBTWPvkSt91jH10lj3qZ2OXzm/iXzXOuR16Z
DeHmjuXLKCxJZ6QcsCIzM5DaD8X1x0Q4BE97sl59S/jUqVM0ZtW2Im6K/kE/gMld
AAtMqEnugVJSXzpOy/Xp2SXcCeO2AAJ6WW2XrFetCyMr04q3AjcJV6h1uU/fDsd/
1oqG7htD74UTv8VJnx82DImAIMaXmufNHS9+8SCj8eGZ+/Uc5fFpqFr5NQWdXt5A
CUrStUC1Iv2SUnRmxqxQw+Okq4GLnXpDTZvZZLanNNuHlhpHM7TU0Uvc6suN/+Y1
DKF4VQc2uS+GfPeLhDijjv971syCysuSamDitk0iM3GBBlZBs5brfULvniDMVm5J
Iit0TLP/0lIluuFOj4K0LboZoo2j9EkSPE0Z2E53ZD3YTaOS1W4K0zdfgbI/H7ib
G8hj01b4gI2gewx5yUhkcMTT7hVPTDRpbgWQQqhlKqWJ0sMLVQkev2+z4x02BWPP
SD4Eo0fbN4bcvQOsuJHTAVzpPa6FTZl+4edYv/l8pmCC15FnmpHNwH2zQPgQUi77
vWhHgFVomJEiHrIti9IPZ0H2xnogqjlaitxpowA4Bma2fcYWU8K8UhrTY2ssVjrt
bpiKCCyFL2aqFpR9fwWHiuCKNLHAG/MLtE83QMVnuxZXVT/ql9obWPzFK7YkjYlX
9C/k/sb2cCaaKYrAvPAWJmsuNu28ZAP9ZowXzqtqnLpzb6jUI7qgwQgAjs29Vy7D
4x7Gliy8lz88v76IGNktUE86A5EOmreR8Apk2PxVdh7CN1Amn+4GP214NTGVP/Gz
jEgf/3gzorc36zkGTMkkxkdHvVW8sInB0Zxuxs7P804gphA8oQxUg1L4hF5HGOAt
lUrj1N9lv4HtTW50lqq/CkgwqAy5kiKr0OnVzDnnZOIFkEmvea8d4uEwoaLwXsUP
cKa+erUi4XQ6eB6LplVOXQ6V4xarIYrB1+qmF54OzVc5dp0vNKMVQfC5+nuwoafP
+QpgW9mPM2i05AqTfJ/HckkghyLG75XM8gGAuPkzIxNh8wtj9axC9QrvkHypPfYF
mFhaEm+/CdXLyGYTsedKRcftvKLyf0MwbuGGbFT5dg6sSz3hsGDaQkNj0WKN2/Rd
tldUbZAwLgTWhj9C4LYKxlZOFbYrbZP8900/KG+xug0r494YEr7wsygqAGGIDkLR
X5bkDDaJzsEICgUGea+m4X2iR2O0qnhGt8XgHB50jp5j037BLzrmgv44AoRRUtZI
xNucm6StGkdeXHIStu2s/2PKDH08xY5EOs1r6NuL3PuE+fwopABF3j/9gIPdx4G+
zhJ8+V+H0mi8h3LbRQ2r8HoyaPfNRwLuNa24L3GFBYP6GucDbY2ojmj6k9124FGt
PuF0uUb3yhLo5BU3nwAEsCnDhf0J8FEF8jib9TZbuXokcEbwEmt6rajO7mc+Mkig
l2WzOvZfinLqGJDJNUTA+qtM7c+rdTESdwnqxM2CU1Y7hxRWlD2rPafWvUGbPiG3
nTcTrS7JmNXATeWXO973MhgOZOkmVTVMMWdZxC8sZVasuo3jW2uNpmIEwPBihD5H
XI8HgVIhbD2ZDLr9PmPr+uLl9QNz6FLFoK4D09hAdlYP5yQyn7j7CHKncuN1pJRS
l4fyckZixVV2h4ZMT6xdGGg1fkyWtPQHBnqUg8tDE8HlBLt8re34+YNYDEcXnWXX
tvB1eSplefboogBe/F21Hf48JhRwj0ODJHBXpUGMuLd+4C4EmHI/9GyRHBjw8WPl
ae9yWBu7WM58DYc0PZDEPvbWYG2GK34gIXP8eXV/jdgOnHPV4nePfJiRUfhEUsTo
xQlpI15pzliepZgxONuBtUBVqWwEPBSh+eAYXZ+4oHTKvTDtG0Zdus7UaEEE47QQ
BEg3c91/LA66P3lfWRLKBQLEGsUFSZPADZaY9t6+CDvUSTx1QVZndXiWZx85JH7S
WZ7JLbTnO24ouT35wily5uII6cl4cW1hyJ9TWk/Akq3dIkxetyWIutElwMXxASul
P8wsdsfXp+fns9Xy6yhce63sf++CwGwF5IEBiyjqB+lUeVOoo9cZMeJ4y3DNdfjh
rCdlHGrlxSPNMbIbvVriXBXEfm351pb7P5TMvuGwSTuDaagNQ/a3vfsUx/9uqe7a
i5ZCxX9qyL6Q1CRDy0ybWbVfF9dpLZu3Y86i5wFSQQfIwFIRUnagrd6hkcKnU7YY
NIdSfTgU+4sLBx3A3wbyQeWERPoctK59Wl+LG1zpWp1oEWKDURphWZfzDIpz4I63
4Ps0uAWTH0to/1kfcMqpXc5qn90UzZNaMWMvpoAJ2yN5R5DWRnzr3nGk0SQ/1WZB
SnXU6v3nzuBEQGUG7G7Sc7nfYDqs9eT0GK+pN8zYBaknAOw3/v7r51hij1trJ+61
H21GZzjmwtbmrHsdGFmJzC6z74MXfJT9w7iwtV4Es9MM3oCE3XH6hih4ElsEpOYE
37NgqfeLfyyjg4ZF3pc1BgIkQbg8UGbPVSJMPU0jU+P3SVO89dtQYexOHtqxktbw
ld9vcHvbhuyXObQWW9SwLw14Rbhp5WasLCtnoTAskc+zaAdHktFuH/xGhxSMtd5g
mJ0S0o8W1fRQ/x/6h6oapcwiToqHqvhUixfzQNVLzvYi58VzIIgyNXGdDMMFeQv4
VG49DY/4zLegO9/H6ixJYpBMNkbuqWQKIkXcGtLL5oGt+M7fGuBVkONSCQmFQJuq
VWUlcId0pYWV+jA1m+LFzmmAxMNDYPROZMZHC+KR2xcfUdhwWIRwT78bBtg9/S+i
DPrlxYKIC7OZ3Xx6J+aUEKXHHa0c7OZ/K1FOn00TB9LfmQd3D7+gLF6M53Q03dsW
9K0Hn6ciWQa5c4EO+43yNQUzHWFMoxc60Fh4IE4P1eXhwM4KE89UC6W5PER8OVSz
KZzQOU8E91LcNwq9aBS0wTIILVr2ySJRsUxK7+A7sHSPWV2wzJFNQzVrzClXb6VS
9TOZBJvaqM3lV9s8C8RN9AkvgbbH9uL2cdSfPG1eOWfFRe6IeQ4UstUttFEOMhVF
vgln1c22BUhRyur5UKRZprdXJs0+s1Oe/0GURu7uqh+KCkxXND75SbCjtZ4NJ/x7
J9lftCTocytLKoSTfWvIJF7WZzo8n4I6BUSwaV93UIxXf5ycMpoSljRw11GheP3g
QdkqEAqt7RUVrRFSBgDZQYkXvBr2eQNuQiG9wNSIdHH9qHAcog2uUqlDdsSWoCC2
WrON2zv6OmCZ7gwEr1g2nIt6s0NqTaVQGeJDWEAhb1nzYaYmaGJonwgdru00DXHg
QnnwL/RKoJ9M2dB/PxLrrxSoGRmsAXVmS9k7Hc1cAsNsoZ7C7hSZnvAgXA1X847D
xYDoa1xQ7NCmc8ErDOHstTSxeGYdODnW3AFm0GU+GC3uFyrzg8c0fTcyG/fKy8KI
7g858sGXIGR+Qe3eXuH9fXStl0s4P5G24l5XsQB7maUSnBVD4iPGNahvSU46ATeU
8pFRfr/yy5W/bkLTd9g+6vFSKUvUU5kEsCu7HxwDKVaiBv9p30MqX5F4dMUj1mlT
Kzgtvto1n29KoQlyoZXbkKL0wkG9Ru9IakZkUBk6B8ToM3eYToDsD3ZAHANh+09J
NDMKsiwNwid3Ob8imkVAhJQQK8MfAD1FifRMDEwMm3lfhuAzcfw/pT4/m1/bBqoy
7r0wqB/ZKcx6LQYAFl+9XeVnuhWIOr+rcdkt33gTWqlKLsQfyj1Qte1qldTKe1s2
zGOXoD2N9RQcPiEtZqesUPXZBfbOZEOQYg+eUYGF6xo7mhr9VWJd4HWpVrlH8nZ0
JU4w11TjZHvgmyNsy9ll+x26fsKRtoIpSiZIeSLykG0c7/HgN2SgXYU11va7bzBE
Rs8oh7sQmUP4QjmYjWZN2QMCzGsWY4ToTdDHWFXo/HsUOsvSpMwnwA2T7XmBVpNo
yPoVZnzraPGx2Iujij+erns+EDDqakMTQOXtS7vg0M0U2dqfzWVARR7gjnrQ2/vF
DeJSrXmr8VuaOgubDVmYCVRp6Vvb9UltwPuTvel2TSkJUE+o6foB/SoU+4Md0dd8
IpktmyGFgtk9cc1/mts+OeFfVC+Oj+bOOEaldTuoVU3tM63RyMh+zG5gJdHWilEx
Ok9QmKE1jDrxSw9RSJMNYGLVf7VDfbp2A6ZK9dbtjRtqql19XaHlFx79tFkDm/qP
lMmITWmNxkbI603+HnBrKY4cqXtw1oU04L+Xm0bO+uLPY4sHAUMbaanQOy8OZfxS
tf0de/F5RFnonl1i9jCRzEAIt8s/lSfiHYPsKSFyEjjA7UVZMpVWSOeNAOYk9O9B
xjJMO2E59OLKmrHE7D/oyWH395G840YOeApB4ZbH7/evR4utOSzMka9D5lo6Wn/x
gM5j7RYfN9BmHHaNtEfNe/lhGrkODrc2j8U7c6S5CfO1z7KqhyweoOSh2jYyTFIr
xiIV08Q/syrhqly+Dn32PBqktyom7nJrz8Jrq1LMfGJW4yHpcJp+p1vjXZmeuUK1
P4cDZa7pv1Zdrjynn3JOLGxWLZiSHNsLwiVr4gli708nLAAM/B7OtoajcEyHIZUB
I9u05y3t7KLHTvKU94fpJ2FLuJ5AOYdWdvSCCY6Fc7H08vkdwk1bZh8kFc2E1fpm
G5rrrWxgCkC28dUMG2EOlKXwlUOtgzir4IMmuUqExvNEIDtJMTTMGXcH9M6xI5BS
hYQxj9qKi9TG6sgExWCh/VTzmeY9j7SLW5YvEf+Y0g3GkKnMMMnHB0ej7L19YXHo
tIbTwGQRCRmvY5vIUy7m/J1dp5mWhwCbM/o/Jazv547hNFdvz4X+i5RqbNspEDch
ozfx5yMIgui9jEVmUnPHJdnWVdHTimfCv809Y9yN/xr69O9wMg+Eej6DXhzY08YJ
zQpatFbYaN19VmGldlXMoZbRORtctVuMS/+b+ErTU4LimKqqMfQD8aO1j7BAbExu
q6EvFrs7yRtrJ7Mp087ULvvtffpWB1aUF95g4mTs9F30u2QhNDsd8OPbbTdGZfzs
mV7gghD1bWkvJoutz0Nwo6/Gp0HJ/9yktAPxEsp0tpOyi0cnM9Z68WyOkj/Hx/dr
IjWldQGKyP3IDrzBWArbj0qI66102iU9OOuT2BAdQ/A0Q9d0LYR3inR3rqXmHlu/
Zw/u5PXgv7lZlh3uSyntx6Fg659rryshFICXjFCgM8EMGKl17cjnit5T9f/ygWT/
SvziDOkA2Zd6w4/C4nbbBs4RdPVPcTqFJ1fkNVq2eeRDAa5cP4hM0fEbcGDgvIit
ABO8HnWjw+mqsaPigvOw2OfWJD92JJteboseiv8zozMgUBt9GV+cW/6MSppVtcpc
SoQV7mLi6+JRWMb93Cuv0WLJcEXyRSCPlY0TnAtihyZv+wKGuhV6J/Xz1xoF5FKW
KD71bELV0FNKGkgQ0+TCNkTHJm8PVVlM/0crHIt0mYoE9s22aH4VXtj2hwNFbOqD
lHccrNM6GSLcNiyD+LVkBsuai93WeoKDpt+rKashHO95KkNmsYBLfM6ZtNqwCXRS
TDfL+qEK3TUbQh+yB3Lt31CulXOWBTS5+yyVM5y7Oh2V0IBLHwM2mOsme/2YpU+K
uYhKXOuoZVM0PSK6mNZkWyJ8bqHfWmVk1ibI+1L77ZolzfqJXwl4O74EhV351tR8
FVIBxWseSxQYUb4zwyFGT6hSngPhqqwXlmx3RFN8nqmRjNFX86WSjtiGLle0grfe
wF069ceEuZWxpBZ9KXefg7DrZbv/tOVW4y3Kvdm51uXxKynkvYhvm0f81iRLsk7b
e9ZTzsm1H2HZlTifwLVpiqWqbeNNrQlQdImX+M89qs3J4ep9IeZtxMVgCj+HquZn
uAK72h0T/3gb9waMrH6XyzHlRb4UyOLT7qcutxyx6dpHNC02tGAzUNfnymsdyIGD
TsSTMCv0Jk9vqpvJEJvRP+iXtYdWdjUyGJIs8nWnFDPPwIEf55KRl/dERXu1+JUV
sXjMzpZ24sebE88WN0vDD7TS3TiXsoqDQzVKqjvpMB0N2rCtVZ75Wz3XxcxhYTxo
nXTU4hGVji0JuxhAvNKvhGI0UnW+DffOXaG+AuDr1wAIktMdYKZjS1HEJ9KCaWHJ
wGO2ModwbBCug1gtgMAtGs6r4YJ/+Wkuhxb/wa5rrslf1ZQdbRGVSgUphW53DF5L
vSWJq5kG5W3R3g8pGG5SOm33nNF+idFbuSk9vZWXNWfmLHSh4T1aQoBJEeQ2jzBW
EH9j5UAWx/ErwKRnmAtrBxY96b6vPs/cbYGjCFXVv2ligZR9bl0vZ7Fl756Xpuyo
3fXSZseEZsLjupu5wLhNCFX0dK2lIWVd3439fQwezD8IQnBHu8im8LqFpeiVbdc3
l85+t/6UPb9eH5KdzrDqbkmvkXSbSstZtDi9z1UGabJ3XvGg14ohvpekj0mjO6sD
YT4u/D5cNgpuw9DhoQPSynLpbVJzf62Y1AuiPme7YXgJwI5lKqWLnFEzhCSALmGG
RO7OVQ4JZJop3G4mofESSiFXaMATgLHxN2LxmYlk1SiojgaFTVeETcvF9aL75OKZ
/B2sLXN+2lPTBgL7BV5F25Kr+8gY7WX1k5GqNrLg8nn2RthZHzgxAkpJMXxeaLcG
VZqUTv2NH0KQ7jwMDDfDEvcqoDwROMd5qYyU2lYg53X+ydNhf1cgw5RqzAbl1lJC
9j0Oblh7aZGCW/yDQPv+zN/rzcsnOPEZ704OLg3aDlx0k55qBYQr1a/QExmYVqIT
clatUF2SsNb2bIh8rEHhxImDGpleDCWE3l+xEocJ1znJYcgz4wmO3EGuR7VlKFp8
tjJn2VJccKS1Q3ERF6O24Ft5tfPECmv6Vk/BeZFSAuFi8H2Mp8/7+EPz+3YeVt5d
+KNuZbLXh2YKKc2RVvGaZVZv87sGveTfGJlepTi8sURPLbHX210wZL1CCwYc5T7V
2+UIq0qWPiFB7o3gCj9Al8KEi6FgjJ19Z+0A2v0Q95DA4dg+QBuTRI/xtpFjMove
4cpP+qDoDooJQdPo1uoHDb0Z4LhxcyL0ZeaFPZaWKpEuC5aDhbXEHKhsWtwLk19J
LXaxoaQxHM3gQTlPw5/Ns/2aYk24/WNW0QH/NhRXRIyNAEg0JPwv7oE7WOuFtKRR
CakxyGwXVKU7/jMgqnUU2TkjvxAzaA1mboZEiVQj+Bl1zxkb9EFnFahXTVFWUV6N
eBkVhLbKhsHnQIFIVuK+x4f9n1nHa0p482EzJ02LAXEgRq72zN3x76TdKoSs7+dL
Wmv0hoXd7A8V0aLTNvP+vXHkBnPyegJuJemHf30gzBQ0Ca6A6WdHvMxfVLCf6Bbz
p+a3tXYbboU+A2J8XNXqtp8e5leyJb9RmbdHBZCXXsJQAvx4URQ2Z0z1SA4PfDGU
MSvTWsIdldLXe3s3iH7SqW4F6T/8vc/wSwQdIjj2OmbECpVuKG68YQeqrjk4jGzo
jRPEqMCkwDTS30gYi6++Cpwq+V6Ru2Pp3I0BAQLT019EdbzqVElcqGPXMDYCLGkk
NUeJc++Oiz0cw3rRhrtyLd0XvgzYsdN8t8Ln+KiBsgufZF1Ii5CxpxxWxmywQ+WC
wTzAW6mz/9ZzLrpyWhzGnjWnfCTnn4FT34wy1toVxa2u+S6AIFvNcPRBgfu++C5p
zxtYuA5FiqVylX0k0wP43GKr3hFGCdR5ay3X3XSI61BUBD1Nau6f4Wwk9XabXW5w
s382A5AOw/gDayn1+RX4IQRzhrfdGWtHclGH9+Odg8wxs2e7eQ0EvEHgr1+WiiB8
tO97N6BWwwcTnPE3GRb+GjhuBldod7CaaJ+LiR6TbrVmkN4EoeecoCTPmQLCipI8
T7R1cs2XEY2dWg0ZnfUbW2UO9Ww98dWJ7w3sQGX5oDR8Jt6UmYr73VCcS5+zMMMu
WfKQ1vJ3YzC9hY6zrdn/Oh8BgYixcPegnsoaH9tL/W9b9LaGN40z8uVgCd4Z14jf
K+f6wDMLkEoheyJ7jWzV6gLfCIDZVvUDsvZ/xF8Qjrl0bwrbzZkk//pdlS7l8lZN
DJBn1YiHlUFU5TpUPTTXsfKWq0t7sbQKCTywnOSUL+b89hwXWfugj3MMWDebopDe
vmoHk5bZEPuWqIjWrfvW6pckgs5iv/T5iEGIfT32L/liTxXOilA7DeJFZK4iwKEN
PUc/SVfTdp4+eVSkceDtHqjQenVbbsqbkkRS18C2+OoKvnhRtk0fhKdm+3XtaeUo
kAFBjfaNRPLtbtfQpdw/d9gbyDJHOQYN58CVQU4tofKoLRrgHvD9B6lQCJYILo1G
5+yXCIaE64AaMMG5L6AXHj26Ky/Zh+4s3PwmYrmqL+JGct6A+DCilyA9mF13erqb
0IqRpR5S1hgjaX9fO/ER6IqwN27ad0phgYuzSjwYFzcbWi9JfoEzT4vLjUnFF/Wu
XaMjtf7Uzq8Mfdyx9FIbIpuQ0s6rnZYXUyScb3aS5cBhoJN2Yxbuuow+1L74kgLP
qs4xRDSdpEwdZYCaSETBVP3QaWQAI3K0lQEls1e95UDrbH8GSyIUcc53zHsWS1A8
gw4COwfysZv0ErECIGsjZI59Lul3yzAGHXRx/YFSZPvN67dpg7Aruet/E2Wwj8ti
ie7dbIfdoRuzAHIWCvQpSt5alvqu+Q/6kz5vGKthb9nZzzwLwTOvoC5a4JoKcjWm
RtwRMIl10261IIm06tBHjA6/xLYz25Bwg7fwaCxsXuXHZn97hOGIefE1dNgU1CG6
dQncvLl+rh0Z8l6HIWC3CEcrkPXWVS2ovz9jMbBSQ5OqqgaPC5nD6ktYDO5FGvky
RHKbp2T3TueTXeEQXghHT2+bUIBzZE4CxEHeDaMbWM85M5NuNmK6KuREEagvkCAL
UEsGHXGm/jJLE5Rr6pFfMGoi4VfzXxnaEgDLbQ/3Fo0btvB4SvK55ncLjVKZAsnm
6P8QnqFzw2M0e5iyNIIgS6HOZzPCSivay7d7d61RhFC4InExMoJoDZObLyfy/9Jq
vgeQjWyLBNjgp9XQNF8nnfC9jpVWJp/MleUH42YXuJvVrBVjCyK2dK89Xw6lMn4p
EZ8WRIqsTXM4OwDAYYHqdDLWEUGf6Jvem9/fTYJVypQIUoSj1jqqJe1P0mKhK3mD
2EGXo/bvJEPQifDrAY5FDU7MpZUzUzGkqWDygGDcchWLXje3hGNw7XSOfIojQ5MD
ePg47iHFpWFQpesGlqT8Px3S61eBpsiVKQdNJ4r4Z4XmEvizBXKWvx+dvbm0YY+2
ZT5aLXaOH0Guk+1SFChoWcuByz/4ncNRehT9rQzajV/8ojPYJYpAnx6Zhz53tQLO
+8VCH3GTUqdcBt5GXQretGQGR7ihd1FnPtXu/fRiRbU6mQ963J0CsnQ3nIp3jGla
KK7aba0Z57xTsEKmrN/NfWkXy9BMR2OYz+ZXoDgb/b1u0//Nm8euoRF8kctEXRIo
1IJzOwcpXIKDkAuiuZJ9nnnvuK2RlRNgr7rucxRdL4hkpYnLZekb0pCQVWrokGnJ
aNgh35iPaXBirAT6RtvmKhACpHnVinSBrcV6BOVxyStWG7exSX4hZgNt0Nc2HYei
9ujYF9XzISILYhFb7o2nIFTOp6ZoJ8VwXjKWVuwS30RjGN3RaWU8NXd6rLpVAlVo
uDZIz69LCHN6p715bYSv0F1lwzHSS93JLX9SNeVCnfUwa6y4QP4KzQ0wBq9aVucn
JCPdca+7JldMa/ixKcmgJG5XZMOT3iYGubAvUwalJhuYjEfPuqUEbZPAllt9lyqt
pwPGtQRmaFZKFDAL0tmtQhjtXaQ1Njm+3N7VP8ohfyXjWNYtXJyR8oZqUJ9OjZr9
KJZ/Kg1zWUek8G9g/+qnIbyhx0sM/ychSA6f6Cg1ys57NlY4ishufRaAyeMKpceD
f/8VnwmqZhUngfgOfLzPF8wmpQCOkCS1u877vBw0OBQslOCWV4QJwbDB0xf4dfv5
sGtGZtTBsJpmDyiEQltR75SKzwEMSr/3Aca/BB6PBWPDdeQKRiztl0VG7HIhllO4
p4HbNwcnJhpuYTLZqSH80Mn7HzOw0F3DwLYpMJfbR7UzN5Wy5zzP8cXNV5lgIFem
JWnxyfwRUfS5oydxrlDmxQaRDDIphRY5xNVH4zJ66MeAnrYz1J91CX5tvSYlb8mU
nMrTZRDzxoz9ZQ+ZdYbj6/7aa7yfGp2+UahHzsggIxhbRwYBDOvIkC65OcR+2oGv
tJDPiGnawioQwzs5TmuOO9fX/SAHKt+079ze7r3w/sbRHN23f8Gvp/z0ZRR3fwBW
ujowWTnYIP8j+jNnHsXgo2V3CBKTi8QNt3cVl02WW9htu2rAv5bFER2IPTubxVlR
Crg4RJYn2vkAW/XAUc1tijT1TNaKxsS6yFgstVQs3x0jeuJI3mS4Nn2tK1dFRutY
Y9sQKWwvOhAO2enkL7Vl2IwfI5b98fXsHXYvhf91U1WS7cctAM/ymrUlDeMM8hUl
/76Z11KP2LDuQ2XGtFDlNUU9T8jxmsjvxMa0wU+0On1suqb+P9CfQgUKhs63IF3l
3tcWtfIrbAUpz2JGiS2Zud4F3mXBNIw6F5oW6YgDVN+ZgoyzEK4tV7zydaTEh56D
9crxHziY6XGHTdzqfqzb6iSCDfA8undYcyVPzevXzdNrUEN84R27bZRiZisY714q
9wrN1lIy7OuJtVQxzvQWGNfHCpblyF0k6fl0juwpz5q4kvOBHeMmdL7fIw4NSG9o
TFsyn/CUOm1kLb8qgMJ5TbY5UOfA0GkuYUpNRnCjY3ghBYTYJ58UkF79xMvn8Kxy
GfDOwLDK/yR0+N7Dhg0KjT1fnelu9Xsdm9yrRFbNPnArZIHRdsXBrFu7u9B4sQVJ
trBWzt1PFtqreAdOu7a4cscxvVaX0VTdxyaRAwldlKnPznTnSNBevG7IIn8wraoT
Kl/YlJwbXSkjPuM0AxFMFO/DOTFg8f+NQJPHe7KGw7VW4HbOgxvrowD32ls2uIlc
GWAsG5vyAJPJAQUjpyxhFXUtCQULdGURXMbKBm0HoJAqKU3Rh8rSlw16GBGu0ABO
pISyaXf7gjY+15W/bE9UagL0IS8/e2cIYQyADM1yEVywplpE6z3rlbC/Z4DlxsEi
a+S8eOxmO0DsbMVfV4G7zjg3LJD0ymSiHuuWK4roPwfChGbV7xBJuydkEnqDi9gD
Xu7aQts3PJhK28WS1vpALjWXM2YORxs1LBrj1CjwjdhHNdMYdNkEVkv50bnRj+AR
8WVaSlglou2rYR/v5rVHh0lEbfvmUpp6UyIKYGatf1rJ4Ot82pwd1M2Rqmt/YERQ
EgkzcqsO7AbCnKViLSzXMYp6hqZjJ1cGt0EnsiHCNfoAdYBpYXBwcote/IPwy63p
X8ICaZwtIEAQj4M8KQIQRFSfPgqSlk1741Cl+csWhCwAiNKLQa5pjeJvIGW0Mu3M
hheEt5MuoQHYk0+4/jdaF912pDUGZ5v2rkpv845ZE0rrGdqhHF8ne5VZ17vGOi5z
yHRU52oIg3yIWLCGmhN4XMhuxFNXefn/iQ7icZU6fYD+HwjkOwr7MphLOuPsPZYR
2mkhqA38+LQV+DWUSxG7wlelUpWR2DXa4oMzMzFdfieHimuJnwG9ORXOWTIA4N/5
L3c04PJSNRFrxxQoILWHt8wATnJwOhVejWmh47nwO4JuOc3Qq7lv3wpROiN0QC8g
SzTHLZYeRRmcwFoFWcV7N9JGfcDlygPB5cefauYYtZn5A+8nYYj+MoKcjn/IB0qV
691ilctMMmib8MbGrnslVd4+lgocve2f1bTqdp9vHqMQ5oc6GCzehcm5PKlDdV3J
8eYxaKs0bhe1h+oeugKON6LA37AtAtgZpJYkrmJOzSGB4DNwtXtg4NEYmeGpERDX
D7Aa9561w5UzKNQKTd5gdEpSGtZykVBSLgrwqGjShkjg22yzWiHi9bOpATlB+74r
GmXVnzlA/fglIHyGgCA/woiSkUZ1ztIFWvE/pRJG3EG8XrHeG3BcUtL91W+3QZ8U
Y2aze7FM/kNanIb1MUvjOxJFAVGS99td1rC8n+OL2RTYxmb1GpweZuCJspSR3Lp5
RzTbSZpse3CMveABJV834/I0kbZrmBy3V4pMFd+LG+mLqqdXVtkH9BeqXABvhKWw
8HXV370gblJikwRULjGG6OXzdHyUJrqW2TL1DedUldP1wwDlQ52aZszOiOFSNp6S
6PT7TqHXruaieUeKpDAlqZnvZ7LIG63UIEkN7tQzbVTausoIwLn6txJ1fMC+gvGf
VhjKd8ZbT5Fh4yiE8WRD8SzfjrBnjkUtRGBUHNGvb2Ooe9Wb4b4SUhT+M8XdA/Nj
LXRZVKHpyfyC7ORrsB8BBslBPOd21vtvIF0WY0GMwyxQsDkWqCwLSsnSZdnmuxA3
Y2lm8zLhl2OVDxW+io5GDdOY8WJlTuQEZnEhSJzGKHJ0c8H0BgmlkPhGPXCcoiOL
If7vM/iV4Iao8aE1u2nCSnJBAAN6lg8prro+tFg8kPmoUilpbbzO5KSza/gPBxjl
I/W/lxrSwKFS9dnRkmTaMHT4190HA/W6h7OSN2YHANKdgCDX+dB2JJqOXpCe9g0Y
DQDDoeSMF6OqwUTCSGh6/28bANIiwdwFU2sdzmOXDc7aWiTxkO6l3Oqma0iwhEmD
k4OBgvZ7m4nQnmPETjW1tjIiOBGTC1WC4+5U0fWgrvNb+v3IAALBQGCzN7tftShz
rUgbUOImaUMWYW00bqatt46jdVNningocgqDydQvyYaclG3v8TEAwxI+BEOXVime
N4cGnjffA7gzr6sdFeWNIrzvpavJGTY79Y4ZstHADV/HQwqWvW89bKx3Wx+KLTUl
xuZYCI3JRo1K8CBxTfgEWsolU/Uu8EV540M9EEm1IdjZd45gkb95gbi98K4t/IMp
rZrLd1hEx39dQGbPwJB0zXymIUXGgQFmnGuybg5jSdcm+y1jII8nAGG69AtsDX8v
q0sfQEMV7d8QneilSXEeqoh4v7kP00zPlEHYXLU06fq4h6vCeHKU8rlCXjqNyEfZ
NE1n5lOvT/riHbMw3iWjssMBF3INgxIYaFshfkifTj1fm1J7KzuR5ErbRuIU5uSq
VxB1wPF2xi1lAlODHWXjEVBQdjfrPHtyG7vFK+hR1Ocyfv1O5AASwsDCJZbhm2Al
zyyS1MrDRS0Tdi/pG4rCpHUSANxRXgX+VnkUh/jXtduEKr53TLLbOdYkooM8w4XI
GduazjeQzDPsKCD6VPrYHv1MjG8BnnCxcHHpyACkLm0SRh3YJVU1I+BNIsFb8UWt
pTn0wPLu5yS4rcH/Cn5BfAf7dDolMfqvcVk1Jvu9X6Ffq5tqgMk2ZRAca2TWGX3X
Bt4hWKfcKmGNxC+DP9QXRrLIaKWL7bAbF0F7rc5ZXeV6/JLANuFDdSfeQ7/BOR3U
m8nhDR8HkBK8+PMqLqj8TYeNjWjiMMUFZYiEW+1Vo+EnIsj/amKDBAWz1KNQD2A7
o1krV7vVk2kJ46cmeR4/BwiAvsb7PSdj7cMxi0NWiJpQyBFRJCEbX5t6fYUKCoHn
g47DzrV9KaTYpjcKf02Zm8GXWetoDt+dA52Cd6qQvvqLei9iBgyXU9kHZhqoEZHt
NxBOptxBnaIQaa9/XTXdpj6qoy6zXXdiD7AFo9GaCdFy3HA+DzwlN3b6QABiyTQM
2GHMN4YEQEMYpIHqD7QTk90x4uGTC4Aiy7/xAT2dsYixHA6J/D5sdXYXxZ62goMi
PZDivuTTCYO+YT9e2SrAgpIrPWOGxFgPpjHC7FKEF1oNbRId1BJynlnLULQOouL4
EU373I5Yy94Ywlz+K5tezWf4Vjkf/8fKfPy7tfJcKqyzOIEnUSobhtVeH7qPFw2w
jPscWWa5m+Ywhodaw1Zjbqwv3qkxjyqfaTKJ1gF4Abx41SPl5ZX9kVWr/BRu0lyA
k3dNH9VAZAfjheU0tTX2So8A/RU+h6PLHt4cGXrDJsGJwWRM/i77MFRzs/PHhFnY
AcfNajkzajwRrZp8TWEhXKdL7o34ITg1m115HzfOrE4pVfyCU+V8pa1BxO0ocN8X
CCh7c5LPvBu8wErKSGMaQdSsaECU+gz9asC8TaCJKIQAHoWm7O7KhQEXcy9prilK
GmUEWUT6WGPUs+xG8sVh+7pEbiW1mJU/Nxr6Q+EJsByIMMNMADBFdYVWePUoAtnt
YZc3Zm3vIgjoM/4dBEHQ2PdXZzeoRkz+G0MIiunL3xw4sIiJb8RtiJIyaWIRL/+H
Bd93zWQXQvgUATxgIdkMEyRDHTx7eG10qtCauqwX9b5jY7J+NkXRl55ZKu+exi3N
HaoyyOzbm9cj1xYMUWkB07+dWVQS+IUvyC0rJN6LHhAt7e2TgBQcV8egb3wG759Q
No6BIsRLtC7/WDm+IGdOoBaVu/4ynPspT2c4qRl9+6FsR1l93EqE9ZIGEyfD3/kH
M+UeTWusJGo5m2X8/psnp5s+Xn40bzF5mdoMtVqw5BYcDpPXmMjtuYt2w91utuNk
9WoboqHh3r5C6QMZAyIoKdwB25bU1PeJFvc8ZFyfx62W7DcYES2l8B7zwEoqqaOM
1rOBb2lc94wvvKqlCXuqTdjUXbqZUZY/MOdfvN08pkOKcf9QtN/S0VgXkopcfw8J
gLkkmC5CfoPKDCT38y9Njmjw+OpxN97Auglp4Y2/W6tWGlOfmrvAP/gdWY73eyYe
CeaPDUINzMHM66yPk+Qv7jXpADkIryJAh6OPbYgZlEeuiiePtJy0rGWEm+lnQu6L
9d9fb+jb/RPaEnnTQ81SuOKiAujjd2yrAHFKMLOzIKiCwWPt4JxSRI3QwI2Yc1qA
3xDiOlopmmRw6RCnkrmmFKI/nbr8HBCiS6j4OGAVe2YrjjYAx17+kiLzl9rq/wwJ
8PAt+qso8jLPtQ0tUbUFDIqdjUVwIxpnDk981R2tDUI0RbrGUxnTnB+gta9zj2yZ
M2Ro8DWiMiihU+pvPNj0YCvTRFyKOq+BdkQ87X5iqSgjOhy8ngOlcj0tOgj/3zZp
H+KRM3HFl+h7aKdh8FKWtKKa4dSAPk0RBuH6goWbBG/4laxIihPAGlRfyQOaHSxe
zTWGRgLoqCXgNepM0lASHnogtSjv59nslQM1ZoxgTB1dtSkH+l3BStNhVwFtYWO3
ZOGCFUJs53g7hrgVVSrPxItb1w041xulcBywVjDE9wkxdd8OGqQXcCVvM7hDGLza
AqJSbg+oguL5W+XxLVyk/sxVIzQW7cKzS6sBUmYVuV4mONVZY7IqsT5hTgbegRoE
Rs0Wz7UJupYcRNX75teTykQ4eApagZIPamhIUTU7WGSj8xpo2xbofpt85T46ilH+
2oWfbo2BbB34aEzZPUxi/L2yJeuRC2W+IdGT3nvX/5zS7xSoZAw0Vp5RtznMgKDL
okP+77ObnWKvPvkBoEuweNojAD8R8agTniG6XvgFQI/uCYlqfUd8eRu50xaHT9Y7
BZgGioGmM0rggVvZ7Xz8aq7CVFcWHcoCtQ9IJ4aM8JLQJCQMUYKOAbXZlF5luhEL
So1I/9aTJ6ZWcNUaSjFX9CcHdBoaCAtUfn9aoCqnYG6DrRX4R4JkRd3NO38s9xSM
Z9Kt4nd5rpMdry8O+9jXHSfb05fTcn6RkDQwETY9VkVKhWLme58YhBjA6cm8MdPg
DpeaSI3gYOwN9WTFdJ5RnPmahUdhy6VwPogaPF6ay/vGVZIfKGZ3Z/r1HFk0E1P4
/hUmzG400e8e/DPJJowOvuxIuCoMz+UhXSRiEzQpHFyn28TYJczDigc9+e4jnLek
3EwV1u9g37ZvJFLFSRKkzyBIcGhdwfQ9TjuSdd7gnuJnfWOp3cqfD0F5t+RFIH9Q
a86h4ByCQm+bYH+R+OQOcEWFvBM/WocJYb7Sb97l1/cKGHcqs3DT+FSthiFmvKNE
7d9dAyOAaKQOgiTWW9WWwqWQXvov7D4p7USVI9f19GmfRwj61wegQJKuDFAUDI4s
4nE4MzZ4lODGENs79afSx6bup0MZpgjFlY/IJ9T6y8W6XqKVHNrmsEVs7fepo4Xv
iIWeV4CWqkf1AWZ1C8/xYNyU5dm6pcq9j2nzUGvnWT6sAdCUgLD0f1SAYwg5MiX6
a6Jc8MsKqZLjVqQhC6uWAgu0tzwvyGgWW8lnzWowm82CRTg6soiMfLlkMid0wcFL
KX9YSgKTC+Va2UuR1GEJNl/u9BKxGEMYhbXzgN/1yiMuNUrGDSksi0EPkL/cy1ue
OY9yC3JbeG2VOttuPkRJqqpWrscQUsceSN29/bFeX2qTf/H0k5BWlIv4/0cCpZLZ
YpmF5qGAZFVGVi++GnD+K8i9tzFsOKenEgRYTWZBC5stR+b1LOCCjNcbQlPU8uM8
2lIePPkFNfIOXaU6vmeAx7cUCwPZqGfeP2UBqDLpjAbsJK4SkzWVRLihrNkyn8M4
kaldHJUErZR5AJtQLspsXXYqnLI7SyTSsMIxkwWpJUjT1h5BChNaCIvIA0sIxVtM
kxnZPV3Wi2/N3byPDg9KFvJqVnUXUUCa6F4caH9zOB3mp3mbILz7FgHSTaevNV59
D26RQe/bHYaNAjCkJl46WxMtxoGHafIq1t5LO/bUT9z2om+xXBB5kt1rDSb+ZhJ9
SF9WxwOI5XRJYcgsmn4fCLx6UpzT8+6ohcI++S+4XdrEHxB2TruEviMa5ftmC0sY
nLLFar3F/5wXb5eCEbUsdVLQHebvuvl4Qy0uEHLjLQCzvqOaF/nfXHvpwCt25tjM
68VqHHvtMH9Ag6ozpuDgoPEVH5qHs/zi1QUO7sVh3HBfiKUbKf2okmK6EEfFHybZ
INnbLFeaE0+zyd7EUUHFtzvRVmj18r33I8JD4TkR5DLxjgTyQ1gm6xXH5zk5g8vr
gafvHIjsND4sV08sziNNdY5qr/SmWJfvoMbUrVnGW1WQtIrk7/pKlFz2RW67syaW
St4rpUVKOYN7ezbxTZvslbE7hHZMgAigi4gHtizbgsn01dvNUZ4NA9emxlyJchvf
aa9PWWLionrhXfM643wvrG5y6SJngHLZ9iFtDbWXqvu1rDIyv7oz/iJ57uzROkpK
5aOKuuP9jWBaOV8bpEY+KqxNqkPQA2al8I1PIlFIXbbYyKucG2u5Rr1d9YUT72Rq
jfCB/8awQ9zYklQLCxePcRws/vrhCOoqtcK1mcFvx/WXU2+Jr7dqRz1V9u/Yk8ec
zYm4THrBlpQT6Kc8UpCnD7Q5FQt9YpwBXD1y3+lFdONkj4ylgXr9UzsehSCHzyme
f+KbbDta3zCZKCp3+Xd2kHguKcBl44L2NTZLjfZBIGnvCM8GPe6XQoSLQlbOIo25
vd+paM8i6nIIkSZVwBwjHQpc363qirI7zRaUsIHRTsKXmtze5epKGcHDnPg1zRfE
lhuCEb2cwWOXzZfCgwEm0TzMEWIXaw6208oUOlDedkQzIn0r1KT6p4R4NPpoaVnR
V9D7DRTQIpT7rwLsnXtq+olofqTVqIB7ht4MeKTqHzxuOa/ejTVInm2139m0jHmO
r3jqV72KgfYGnIGz0/mUI9qLL4bs3rGNO8d34UamvkKTtKateKMsp40J0+Bg3O9r
SRCRVy9nvo1r+keEMNfm/nWJFOQlKoKyvDl150vqJ4w4kXgXRJ6O/tn/v/a8XPtR
tU6J5WDrfl1M3X2dU1hSfiTeTa0XqaQ4wkyLhQSc9xVzF/ZIGV6SWGYSR+SfvOWg
WleuhDLNAukSLk+RClI62VOpKs9vVIWD0lR3GRT8nnWVXDaf5TUisajDsDaCnWpK
Cn6Gw92i90KVsfRFfIr2IdTmRCxys3LvMUGHG7VjfXIWSVIlgfFNrBKHoVZZQZGn
aJp8E7xQPXhZHjIVsZIGvPZB+L1lXAzRYfb3hB0vQUoEkr6HjTGoR5upnzsNC2Y/
+e/irK4V0DYn4woVjmKdWb5EmF5iTeLPxpkoohU9/TPo+Wc+STQw6Dymsk7JEI3K
UGD51jhF+Q0sEwIx7+M2sOfSQsdEH0JrO4iLzsld9jm2jmZcmdFwwF2ZUGvAUUEt
EsUx3umY6aacqdbH3RAuOod3XKl2maBUX2/z1CtsNwDugTRk7lzAbaDZAgCTmK4z
tACre2J03jXuxrzoI7G1lCyD7WasqjOfvXJvZCygziO36vQskmLwlmHdE4ThGaEL
+8DSxUC6XtHJE2PZEkRxuEAmPBLQ0lHOuWz1DXwsDjhmZUj4GgDepJez030ffJVM
ergzqiKg3TT2rXxftbepvnmZywLlyrppG+mMFL/8TdqcMGavjIgTw3FhbJhFwzYh
oTJ7tgpM1kE69IxafElizDNOCFWx8D4elU3DqzK4RkVnJz0AFeb4EQYao/ebipPh
hZwP5M6WHD3wrIVEFFWD9OlxqEAz2yPIlPgsyPil2X7jZgwkRceHXJ3RSZ1lg48N
V6aEPjIxExOh9SgxWVodhDDVmzveR8zwKvVKxEO6O5AdpQZHwS+drgaSMOycK5pM
glcELrn8kxQR9Ie5xljCz666xVMXWidbZ8wbuW0UogL+0loXk/8k8X5Qp0RHxr5J
jg+fTPgyA8mFFCPktIHQNlkZW9JprtFwigyafZiVCILwVqZLmPlzMoKv/CeY/Ehv
iTdePy7lFNCZt69BOd2VvfNr57GwTadHrXUfue88xZbgfHKtp9DXHntwggzJrH0A
6ktFBWk5HppbpsEnZODcIU1ixm8XNCXk+S8yf1NoIvdIx3r9c6Z2/NfHX40t85F6
hJB5TqvsYGbOxBc3xH78sYjcZmlgvBEQGZvWfrfd2wFavFQchq5wEHCjJjorI81K
7pTBrQTFyk4t2gb1tkGqKDMXkqn7I+w7VTooX5HbTe08rJgEqnmEJzz4RNwtDyse
ybLE5y2FRs5EvguA3yqXgMmpukA7XGA+yAh/iETrcu3bBMPMh6G/q/Q2YIaTfQhZ
vQt7peYx3qFSmWPHuE1J1q3DRzhw5/64bIopmK3ou3EGDfi7M6HNSpilY7oW4SPG
6vpM9Mpiv/K5lcBhNLZSshByQ/9uiMS7nU62kfcqMa2btOoWycj5VlzAjXy5VgAk
+gJVe11DIvjVDvd7hNCGnKf3wVQpcScoddWdrRDqTcr5bRT4cx3vG+a3LcsAbDl2
1nP12cL6sBLd7yK1pBu0HehS0+PxJtvyTSVVFYNkaWtPnApWPM7bEmk6iBkdh0d+
5uGQ8OL9B0oEizDOoaSgC7VdIJZCopNnRTJSbraG3JORPcvnzbPhAI0ZrAiBtSfM
iC4XZ9rfIO7sTGewNQC+wDB/rs7/9Q5OJoTk0GKPfJZRN5o5b0NczaeZeRev6TYf
b+ABApph32DKIVEI2DdquRvLcyGG/rNiwjPpnm1EcyvFOrPzD+C2FURk2U04yEDd
vMEdnzts7hqaiKCBafEPkQqGCTmkr4/A+BhlJdmq7SU3Vdys5Jo5cePQvCzgdc2A
te4rtzWkx5vJ21FxkxzpXqb44DgQzvGTwsRgxZqXDi5WcrgoApjognliGEynxdqm
hEXyIlSTgDmyUQ/wjKDDnY5dyyJvFd2cAwNl0R0XRPwNZdjiF3cbnSYvBqXswM7Q
gc8IKFhSX8znlww0HGifMHlozy79FamF/Lxk2sYfGLMnoJezlDUVBuJm7g84M450
EO049wjmesXflNASYqR8du1ifEmeNL4EThNHADo+7BkHRQNujfcS68shPXY7tiiC
ex87Aq/1DGZoFXwSIOkr66VLqrPWyPO8dO243fH7UNPQGcPBNhrZJuFEmZW+rb0h
/0Asop3wWIrfP48DvLYwXQ4I/H2SzpKUKvcm7QvfDCsQ6hVGF8MXtH5fIYQjbVZQ
56i/fE430sjeemoFOY5Y1of5CVUoa5cm8PMCPdxASpwQxEXlU/RmiOuks52RvSEv
+4kqAx2MXfGHx9nJhsDEYMevI4De3Bh/7rZeCtLwU1q4scwq4g4lVTcktmlZ8FlZ
szuENC5UzqcqaSp3dnmG/OIxjI6PDq7wTwVAoJDKTnU4TvJPUUvjZGwxyeHoTFy6
3/9PTmwTEec7HI1Rl7hewrR0mG7VkQnuKoNKsTQ3FFJRygK0RVu7tT6iaVMgYmGp
zObV+MAq4HgceeZsX7IcdO5vcRQ1/QVMhcNYG9UEYT6p+Bjr2ZHEIDqwQdDpUOyu
NgIM7Ky3EfUMz/5hz9NlwPjQribIloF1VqjKMW4xdc2rx12eANMM7uXDEgHgXe3M
jER+sLayjB1I5eyzTPFbsqzWTKT8HCaE56QQtuHIlxJu8yUGvSrTTTcNPgGGVwJg
BvM27yaHs6OvVO/Oc1tflFzg/+7xi8KQ5M6gnnaSrJgf5tDW3GBO0LsmfX108Lj5
H+QrRTDeBItBB5FcFId0bVMaXBVRWig7KZFDoVVs5sg2/hJoVzk1zUYy/2zXldux
b+JZHSyY6mKldB+biDfQ559fa0TgUISXfNJOo9yY1lDLlHv4LBErgCl6ulS/VtMW
VbWK9iuc1c9Buydos48T2OisNVVd4y7cu5thLk3rZVnjAQelVMJUbGjtPmdc18b/
v1JD2Js9eEt5OtHGjaL8oMoYxESfSTFRSe6X/446leWqYvabaZLATuCq/WoUSV96
U6QY27Vt25NexEAhKRi8aIPJgXjS5hZgG9eiTcrjEgGS73gk9JGfM1r2V+0VA4yQ
manlrU50OCSla+ndWLpJrtBauzAK7xv874ESRtbzlvZr/h4AGnWBhxG6M1j9aGzu
UOQlWqkg98u0FokZ3VNmT/KFUc1XiTwF/eEyrARlay9lftYaKFQrNxJNUDPXbgkz
Lq5VWKi6BBJRUoe5OFvmxw+xS4aGK+K/JwimQh+TI89Ql+fNcU0BI/Hb8VoMZ9pW
JCcMRi5C61+7IfzIg1mdVq4Y4Lzm/ZB+rX1qmrfzqFPoKJMsaXXpYylVhWOmxx1w
XOqjnFLEKSUBDCFSebkv6Qdal4AO7uRubB0dUKSnQkEJNo6N56Uyog8n0js9bFvS
3lXuQiAcXKzYEH7XrH79hvNlBuVT4h4thtZxyDR3rHmpEZwb9LCX6F51SijmKajA
WKBMxvJSXuVwfj0a372Uu9XuTAntc3ES+kwmgPxlHknZIvh/nIOae/DND+09NnG5
DmD5hrrZA1d/YVLtxhwcmozevG0ZgwKSoWPZQQbIOVzRuq3s9KSrZg6xUjkKzEdr
apZfwceX98eZDAWlKXgaphssQtcCkdd5srUOrkI46B45N9UO+qK6qkkdkehzszX1
iS89ZjeJ3Rsgl4Gt7iw+xCfbCHAq6LrVDgH+7hMXpl0NGsjC0FET6sj4wGiJN0R+
zFcdX78rt1xfVrQ/HrqX61UdjKDPF3vLT7AfmB2k5m8b95kjImQ1PCTIrhaTmKrF
U3Xe1zeBXUWddH3+dJ9Bcn9lWHXqSS+wBuYuz82IvSvnTFerQg3po6yCBAwHxnBX
4pPSwcFNrxl0F+rZa8RIb63mYDwMjTRLD+DjZVauaWAJeIhzqt7KoCUlwL1EtLe1
p2/+QWyQU891eHD+jQgD/NJQQMZI2J2/AzbwFYMy5aChYoBpwoG5bsGQY1prdmaj
uLd5b3DA0822hJ6aU+0jZfXsHaKaR9oNZOeqYvTQGxliDH6sX6Niv8NREBdzAt0v
QJcty05SdaZ3yOsgBxfJVz/l94yjTbB1GGLjMoiSl0hONrS70C3q4fqe0VZ45w6s
f9lvRK3ue1k9D4kxQxMjGiD2RfBJ5RRisGIbPtlA1Wgp2Sz5JO0zbY8wR5zQNiQE
LvGdDlzAjdqxfP40/zjHCq3s0vvMVIZhnnCuZ8YZx8Wcq9XD7jrWsdrO/zRocj3V
TFW6OZndfzelUJwDRrDwKJU8ooJIsy/V6BpX+3dC5mfJlQXTRenJpPaR9GjoHa9a
/nzqDTjWvxXwPFTBxK9irLhgj7xnP4yyLhOxIf1ejiCFh43sGkwWa5/caZokTZcv
c9ye8yCeWP6vfrLTJeUrl0GLi4qSy4ikB/+cY80PAwPrB8TY0DOeXyDDMcP8iS82
XiHsium1GZYrAa0TuWH4vg+8eywxURP5tJg+bNit2ut/sHht+9TNVYWYXIsvvjfX
76iDxIzVs44+zU2WhPOn8fvIXc+8mkcJ35dPMYRhTbwS+IA5hJO9aogFH6PCXIZk
SlbddY/IN/3KtabyHtFnT3RhjbdylXBGsOM9sg1GtQlrDlHKD4g1ZVvL6G8kYQWQ
ykvgLfCs0vgRj7rOW93XzI41u4OLlKXE0ccKzdKDZGsxwXm006b+oRES3ePv5Mmv
2ZVaKpFoPQ/6HNUzOftc3SP3UoAuGNDE6BD5zSIwgueTirOlm/zzXmuspCiGgaMy
5YD6h8k5jI8HsZMGic0ekAoXRrvCopwpLkcBfyXqyF8U75V7AxIRAdsVHHiHjyRg
nsU3892PQjEw+QoE6TOIsIaSsBZef3fSCpcmXFbF1HGcNjCBlPHxMXAU8Vf46eo9
7jMWfh6lYQtopUMBTMvEh1eYW4S+y0r4e3/SwgDUeKbjOu9qTdoJstJg2b0rjQ+5
I93VLbldGXReYJ3Cq+QCNAIMaRvfDnnhpdqdJVYcWysKjTXq7/ceLjHmmvuH0ki7
76cfceHcQPRjp+MYXBoTvPflGtgc5ebrtvRA5ArAMHr6TW2voJrqjr8/dVjGMsft
yPS1RVsaNwxSCwtwReADYZgs0wrG321B32rZ/hVhUDl1tduBU0NjfXNcXMZNdwKN
bFTvTM3jxPdXg3gpxxw43CulaD8W1D1DSlGVpoxZerWc7/G1/GManxQ59m6Arcdf
PshU/tWGkX1H5oJ56KjbACGsv3iKTx12JanbaWpXiVYd+jtzARpI2E73P4u+olb3
N34PaOQTGofoI70pZH9bFat39y8TR/l/n91Tdf3FkIJr3tlvYWq0i3k/D/fTPAfa
JEl7m83LoonbypOxsdz9L4JP1In72M7IFk5tHYP+zF6HuHZr+1Ao21kS5K++WCzB
wMhaNlM/Axtd2r+72SAzkDvJLg9Gg6XKpDGaaHkBRAOnrCxTl0kAV+Yt3Lv7qqQS
aF0mVFq4i5s2sXlD3i80Q147r048KIK1OCgT/eCmZx+u0pH5kS/E6tUvWs1wHM4h
kBj2stnyL9p5PaWpFCrbSb0l5TrTP8JE8rF5CVOzfM436vwU4Ru+DzaHCrCJ1eHk
XWAFpwjzpEaLlA1c1UhlwWjTaQieDDTeATkRhzihufOq0k2Yu6/WSjBH7NtJwoq8
mFx6g9Byrfe7JhbOatfRtklmq0MQYzbPqS/7AF7oGm6hZGXXimIZs5dPTV8VXGSj
SKx8K0ANhfcKyl4MUKbUYuxXVq3VNKGkTrm1nhALBdEK7ILOe5tPCrmn1h6gI/pt
0P5YKGanRGjGB5lgMN8+CIQ8+/4wjNwYjYPBq88CV+9P7H2K4WgVzxTmv3UYj9De
lC/xmK3eNk4jfVpm6to+rSqS0QmfqdFCgYgsNWYsjRVZHkUqkWhwpcdMoIO589K+
YTclshmC49rXJU3P/gSm32vIduD+PnfqNWRYkFidYsFVKmJVCmAtvvuXBSZtnvlT
I60zTOvFySGkAYUN02Z2tr8uu31mCXpeJFeXAj8ui9yGzlryOk0TAK77BiOt/2Fs
T4KCZSklIugoZVCqpdW5A83KE/ZyxA/DGCIzOVxzJ7Ah0qziK1913iOWfhWAj0Ph
ZCqVkmxcvgKCKQgHR10Wdsd60wHRTCqEz2Ow+H+A4WLyTYoLKld+QS7orPja+e6k
7+6XApZv5pRDu70tGRRV3MLW+TpWovVP/3Z/2b1L21iAIpz/h0IV5QmrZxNCoydu
+5baXh8kSSVv5lo3b39JscOIu0v3mqP+MAqtuTZ0hNd3DXztjBPeQRaee3nDVxz0
e+9SiQYuMqamXshatTHEWh4hCBN8YIxCwkODBmlVxUqZbhAW57WgoPrvtMcB4U+V
tUF/PeNXRFmyOA52UzHHGp6hpddbDoxKDvXIpmhAjDF/YLcaSxNZvdCAj0M9o0mI
zhkOw5YNpLYQ+dbqYf++oB4hhSOEsKnhe01chmebNCL0P8qMSjmd+9KVJofsXGq5
QFv3/cZ5mL7mBXjb7OpUXDMzdlcpdScSpTGrQ1bXRWz/daW6S4lsktJsLtbqokwV
0UaVmBL0YBv0IxCVhNgQ/ZpD447xg32HvPQaTlMDu8tPmGhVKhYUapLVxemhwy9N
YjCWqGuOSJWjCgk/MEvjLTXSwatAL+0MMyv3XcpLlIIxFn3SV89zaVO9H5MwLr0r
6P8v57rdW5Yf7pNrtGSW6u3IZLRBZ4TID2ygWejfb3SxT8WvBQjPhvEwLyXbWXso
/zObvWsnz/fzIc6eEeG778dpkQFDGonx8hwwgi9AE2Pz4DtMjttaFogKLFb4FreW
5mEezUlsw0srrgL3ZETmqWnk9mvYpdZXUfi+q4y0QIlHrwsUU+HtKV5qce3PnbEX
xXrj5BAbIqwWDU8nI63alxCyAqvHMry+a38JjiE961reLySkoq5NJmbZSpNNbpCV
1P4ot3pB4RP8FB4nB4eN/4iKltJ2he7SFTnnHQILcE9boUB6u+GfmFCYEQd4+63u
MbgeN/BQ59c5r27oVYoJIPN8aEUuaHVmayckBzml7GJc/eOolNyb2TP8/hzcZTym
WJLmYRB/3qInuMQGkPJEMb3iVPDLAP8fMNxUPO1wvRHEs4ZpapLUF2jTY7AG0kfu
0G91hLAmSW18QMbiYLZTfxzv2qg1EsHdIoZEsR9uhZln08HLnJsUybb3HxIOpt14
BqUcgTyMh/P8Wyy5UyP0/WY0CdVrQi1QrDqjtkZb6t9d3VbtPufWhRQwDOSGn21a
ncVORgJeUq/S+xMeYfDgaaQcOQzf8wvWPxt4OAmYhALKi/eWOb+qfzaR9Ha0IXQl
RoFy0YCp93pgcxDpw68fnu05zixYcHmdmxmneJPQ3MoodeHM96SU4IWurjmA/+VE
omSAZOjXjDc9ZfPA+3SQnA8/x8O/fvX3MSWjnSPmzmffj1nHb+kRjXkhejZo2qCq
U/xI+GJIWHTR+syRLYTplQp1qDZpbS0tyVoJ+nIz6M/iCuIJHl3gXr09tywwGML2
Xpgs9SOglfnCLVz3sTnVHcwwDU4dB2xIN4Xt0JqM+SP7NXvNp3qMgg7Wkd6KWJf6
ncM1PbaP/JMgyFCTbUqepmLAQbC/nq8xV92FWGZeqTEWGy+54sHuvn2mgfVKoinY
RruCXXoNfMU47k4ZYtUxNJJ8CfwvFfqyLFDiqz77yhZztzJw8TqFkFQgI1OFn7CX
ct1a72f1c9ocuItHkPT7OXSmIFVMpCikZRMe5lKYHjITxmw79SrmhKrRJqV09KWM
C/BDFdMq5/V+2OrWeLmq1q3ipZ4H+8QPF6Sv9G9V5NcANp1G6RGj8Etcx5RxMiXP
HjTlFonZV8F+aVsC5hRGk4WlqfylKE1WL+JrlO3lA9C2QNTSy8WbrMW+Uxs2VQi9
ldqkzRZztiCGtCTWZZ4kKARBciGNFkU0WXoyKR1M5ZE75gfHKcJL5OGaNRo5FbhG
EesSNGj27Dm0wYtPd3jOTUBGrMc5kU5/G8koaknIjXSxZtxiq8pB1EuvulYbbmx0
zMZl7VJCQezoe45XKs+vT9HW44akm3lVHDOhZilYiuXL/VYI4e044R1cUgwYQhwl
g/wkPlgf0i/yLGckQIT/3ejndZiInVQg2DZD1bliCr3CinN00PV2nSGThS2YYRql
7ozv4gPtn2zZPuMde7VdFRIZAdGw+yN2EkYfAEXnovQUR7+KNc3mSse7/QL5URFg
GCypJLBdAiccj4Rh4ofBzcf2J4TwUYX37e5OI/7V7nKgUYIvMT9IzE+me8uCoQJT
BY5Fojyw4yN33uNBG2E7VKogwy3IYuda2YJCI8YFsoPktUn0a74EFil4Z6/p+RNE
Wmk3tYZ67XUlrG3plZLSmzhjcLAPgmt7Wgsn7SxHSsRV7QPPt3WC6vRn+uWiPENb
kV2I2uLUR3v/KZ1/Zj7A+ChNLQgb8lrcrBovRnPgAZouwPUKAH3+D/NZhp05mwJ1
0gjHBiCymUDeD1EJmNM7XOYgTSWHkq1/76WX6a5ip1KE8LE6/yeO+X+rmLOFzW1R
bR3eQgSV4ar1NTJMil9nlq9TVONtHu0Cj5jQjeGryYIlAmolsSMjyCD0je5OIBZ0
tY4e7h5wCt3q4HKYkugEv/KXTtW7SMTMVKMDneo/KBKHHwljnaQ94r7DJ0r2wHfW
OWQ1JoYxSDHiss2K94571gdzgJpdt3SlJ3yu1IUAUnlI/MgCbOeq0EoHvsyZ3jMQ
Ih28EwncqVCHv0raOiNN0Nsd6L4USq29zVFwf5ioL5L/ROnXuVvC5CIcX1H9bFRQ
s/yBJjgWPhpdJNBfHALXSLqyQ2PCRts8rbAgHd1VTzjudzjUje1vixrwCRoKsOtW
cI/W0bGJUbI4eAl7zTe7uNluB5K9OHsrBDX9TcSUUU4eqwCOrkyvazFQCqP1vg/T
lxJQOf2fJSHU+sFpvFq7sXT32wdAYWgvex243YLrm9trnrcVzyj/96cmiprUPCIp
n0IQhZTrOYxgft/qFtX+DDBARXhswQjDBOJbhOk2kAUN+mfbXPUrqwQk0gnP1WuG
LN6GCHzZfvNdH7jBl1d4miQbld2hEOlVivo+NHzbWAwELNqW1xxHTCalcuyVze+6
DFfN0F1pp8QuY+5t1Z/p1owiXHODJkQCOuLFMq6uf6xGLbf5XMgMf2scm8ZoYSwN
VhZ/r7NVrtj0Sz1UcehVfBKtkQpocksCNTLChKPrcmLlPseWHeF3XjEGagBfyLpc
aKJgTqtG1Bo9RGKODYr0mqdv/ZqDj6+1xfHglo/7dvxEpRaGStHl8qA8wd9qSSUE
GnnKa0szKax/6ocmsH8IGg6FiYo/e1zyFu9XlcD09otIx9ECz+lU3JXatbmFh+ZI
eTaggHztScQVOc3XiiOtp8xIBT2GWefPDC+YmgEdvtnQcDSUbDaiN7/WxV99KsiC
IomLxyHotJjmSXaWQxFsPX7iQXl4p4wLQuFRSdEmaOZf8oqyO+BVJDepZlvw6nDF
UXzP3YMA0dhLgHfgyZH+NP4h822SlEiQBQAkTzMEI/MZhnEj0oDLcwWbeYKPwoiJ
4PPRrtBsyGeI7ilCl7WLjyK/3fBGDRKZezfh4Cz7L50yGPV8GhNk0+y8YvkRLpH9
lkAklWY9nPVDe0P8iTruPgB6I66FGqDk8ypa+OLYU8r79K8R34cK0QesNc1EcXXQ
5D2CAHiDkrDWs0dwL4qtYtS5bUmu7Bn0YAG69WPDQfNPunylIVRgocgBbOprz0NW
217fRVzng0+xHr5ackIBX6Kkb5SIrUXTo0cZb6wMK8d3NHSu6S+Jd/9E46tjyP/o
eOLED2Ypv5xzspJHQIwqKoxBjda7YCBulVZTS7nbLpacOb3Is/uxeLpKVenMtM97
ql0p6xDC3SiIjrYboRAkSUkhwj9H1bfJv+Thi0Kqyma+zGhHUAIp28JoecfaoEnX
2EwncwkY7RZHqOU+OA/lQN+DcztfxsKLWLymBdQut19mXIRT6X+DirSL3bQPAA2s
QaU25JjAZqNoTOLJms3VSdBvQ8QlDElAuI7mk5QJKq6qZdO6ELoop037NUmkXOYx
Dho/FRC8OUWENHyVwnZP5jmltyRuT7xS/pJ2q0KiI9nfICM4E5q4jDGWWdZZB/Pz
axqpRnstkR8FZO6WXBvQdjkbSqOsUE1ajKwC2X0J/ojBJ5BFZW/rUiq0h/qvvckY
cqVo5XanNX0b7sidSJdoTRbUe0aWKekaQkTriuyuhg0xsF4XYkp063xxW4PWFpzt
D7D0tDuATxORi7S3jHL8cbZ8b9xiRZuqCEWW6Pp0n2hnf9k8LT8LMx6vTUT9uNpx
dptlx8TOIuteoAJ6pOS04mzMInaSlnP7vXLpqQ9aAKVHDMfkTE59Ql1WQ/bu+vyQ
AbVJ9gH7emI+lbWybEtBHrCaDBv3YG4ubMp4eVt3rob6+ZgE/EneH9FjlXSuLn4o
bvgIKQQnMH6jfqQnuxB9jJ+2DyvOR2rNQslP19kCwkj+UC54Ezk54ryDpv+UVQ/h
aSDpQmuFns0hYyvv18WSeDX/3SZ4opnuFHEKBn+uUwanLZWlc0v9TnKLvX7ewx8x
9AK4K8RrdJ8Be2mp6CyoJOIAkRoY/Dh/VeaJtwRQPn9zDXIKJ2le/7rUJuuUKwsu
2l0zLydzbtz2JSvouHs3Cqf56XFV81sglko6K2L/KojFeS56icgG/c1q7xFuN4Sd
cnxCO3pq8Gz2jstP9p7/zzpuCSUH363A4w8HbAE4cqeA726JqvZbMZsRZshhJUSg
O6Zgtddfzha395x2yf5GrkhPSg2Ael0R/juuvzasAtpa5mtsaONTfM9B0B6rZAm3
EJoXfJ9SLKe7nBhvWqPV1MtewaK98JTXiGV6bBcvwTCxGpHTFINwT2XUK+KCu1HC
iLN42wQXlRl8vW7wjrTGUJxijHh9HdAc9drDHaiKl21fEKmC4EluPxD/te8yijaO
f2ZB3V+ZYMEJ285VpyufVJs9jGAFXldqP35UaHU5Ocu1lQF2ZhEC/2FcSkjSUK1/
FVD21ulLJE8v2378T1UTFfgY10tQ7DBU0CFJla25uRp/FGEA/8mlCafaEjdDTqZO
igHQaMz+KrZMrJItFlIdMitBBd36NlhdGu9cZHVuRjIju+pP4UoXRWARyPsnOzVC
SMIScubaL5s2jv8g0gOzyRNDhOegllLPDNXf84ZR3DfZqpfZolg8m3GVZaP3QqxJ
uukVuzkXAclIaF4IuBj/+WoXhBDX1J2kDit/dMvwl6hhpOCXHNDMs4DQv1H9xzWR
mH/h4WznZbtLx2OCYz+oiYOqvcy2RA8s0xxcyuCWBcmyMKgHGNKA7Gv8jEVRhdiI
YNHWbHdupe8xtPsnsj1Fw9542sgVLrmJFRNAlZB4/D2nnnE3LkSbSFuxYeigw7jc
RcuPTohiY0hyHjkC89qR5u0zU5s/Lt0N9miN99it9os=
`pragma protect end_protected
