// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:32:02 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Hp7/HcNDdvpOUEq1yog9dTVk4TEk9BuxREXFbtNSScLR9AVkk9cw7C+k1ZQG0Jm5
bhESqMg7/iVmNgANWXzKIaN97zwcPY1o+lkLXKXhzBpTYZm+DgfE7o/bDw8bPYR1
HpatuMMnaweBaoyZam9ZzVA1AfG8S06O0mWNpfxWoCY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10976)
F3dKtEWIOw8141zZCReN9vTEkNxXeVuKyaCYieLVCaGo1tvr9BhWzUZ9505bDwz7
ZM0H6w9aGocFovK38uxaxIJu3olDZOcxTj5zH9FLPdS/6T4sDAl/26LJbC+wwRTe
yV1sE+DYUkaXzelPl3WpBnZqIXH7MOVrDWsNJVuRkGjl8N9yPmJnk31bLYbMA8tu
/FcC2o/fN6JITb1B9x9j+zdkU+Pgj9SsElBzBm0B2+ucK9hyy0iUah04wOa+T48t
kVJarKkI0Vg37c5kC6uaDCWHTdjtizYgtAt5nixmFd5TDeSaPMpKm7udOg0yaSsO
X4bwWUmTmr9RAQBfxtyHP+8iYCLgSa4C2szQtnS8X+dm2p2ULcHT9ppC8bJrikUa
ONQ5JaxwynvS26+iYGDPXI3UZY0XhTVDJturE8Xltna8jR4X8NW/IDxYBvlt5JIH
4M4MBaUzHQKpBtX4wgh3Oawo8CDTlnkUJcTZI3syWe6bLkhAaKQs7U62LYqV6Bqo
yXUuGfVjEdK8TdKbPfqx7YG+Ty8qcCH3qdr4YpoLPoQZXof526XZ9VXZ6XsK7GZ0
m7ru5xpSh5wmi8BW9M3iNn39gNRjyAd4L+1EB68d98uPlMTI+EFv/ED/XnHFqw5O
ejKL5bdGjR+R/+x2rjz5sjaVRNw6RS31l/EdYvgmZxiC1JRQAMjOwJyqsBMtsPms
WSjzM7VnTkb8255GTZIjNU2LNSY8zP+P0yvm5943Iyok8NrZZ1Tw/mIjC/YDMW9V
3vypOyIGehXO+4ZqNqwMq3dQ1LwmorE1MhfvwmzWtRO4B8tnUHyPxfJsYLAAoTeR
EngMj/dHeql+p+I1k45yfmUOA2kOzyjVBuRrQPv/bfYdKVFldh1qT/O2bC0G4SUZ
6JMEYjQhseoUlTvpYPUZf/wcIzRQC2e24PvMmEAkeBMQNJJMdr1CHmmmV1RLFlcS
HYkshvCPUkFylPl2htl4bMJtW/+xH+iEVxP8CA6iVR7VFtK4ChdRe57gx6wR0K/5
uOIf/HdVxBe5LQB3fGFMfc99J0Kre6v602N92uTH6iWTvvc3fn5f0xyJ0oYPIBEo
kacPKmi5KA8NJ9JwWtU/YPCSV5CW7/+59LRo6FLJXvnobEfZpK2aeryyTmpLuQYq
lb9bgdIYokdpa6z3r+gi5NVb5T5WQBUMcbGT5LPUvIQZvRyhqxJmkYCrpgX7jS57
Glm+S3BRuyidViJUw1CKU06O5IceVCQla8Q5S/AXk4CYA54DCX5+r1EIfKFxhkQU
zAAdPxhExmmQASgn7t02OiIpTjVqNq2m6VATqS9n+fayRTXHBX1/pR35rsl4GKOu
9NBl9FjErhPpiTdpRxsiNqsRp9jmIIPQyZBP66HW3z6lu5F5SXbZlnw6SL2C4fJ8
JAfXsg6RLxJQZJG6Q4JaCUzVBswG62pROFSVHI4SnPnJV6V2ObnkWgNy/uqloO33
WWWQLrhIeqnSdSxrAyLacVzp2sDbtIY45utCvpnpGfShF/eHwNsuFbu1h5gWRQWU
AaOwp+p27zSpnRYH7gnMzd8+wHaJdD23b4EwMiqqKiaFNV/7rsvj74H92y8zOWw6
gaRvl7TsuSglPvGg0AsJAav0vwlk8fWxZ66lj8vmXjSSjOzqhIp0g8xFwbSiRscb
fOzMHpGnnNGf+LAtQcd7ciRESiJTdW2roE9v/H6z17JOEVjZoQ/+fkumFPv6gr5Z
OSnLHXNLeG0g6XsJK3zvq3+D7cT8j+H8QuM5HCZ3sqaPtPEe+qU5A3RRMR5Jrnqj
P02ERLvpu53wFvCNAuVInQJriUFbPpov+Jdlc43ctXJtLyCd6ROLjKHy/lGBJ4aH
uo2mlIeNiRXo6w96g09dL+rNLavIAMw/pyDypG/FiJ2B1zSXHqwNYtl7/dUcnh2O
tt3bpjAQfuls3qZVWkEKBzc46wHVrcMssyDLHKBqjDLNtnWB7gmbQofsg0U1UVvu
0Txy7W/6NyUKpeoMpn7FCGYQn+323rfsl3S+RU2bqs0VE0VZrKvf42QvPhdgUZRE
CVUA9kTZVuRmN5nImnZUQq4EGxqm6bVQxKo+TxP/BqSSQt+eBZZ9rSyVEzoFhz0B
XBMTB4TZVbsapLHWx+KIrLGowXa7gJPA8lS3YU5PbLSw895/Wapzo4V0yzbAelj4
0BOTIInRldewey2z7vI+0W1wf+Sbu/8EsR9AWqD7uLNgWR6FTKb9CwTOE7f7GU99
dEfiRA8jO9/GOe9wBIHPSZnmUbnszKbAPTUQ/IW3fJOowXA1PQRBcJTjwS9/2mcV
jt87UAeW+1eeFkNFbe9LlCcbQSSi5a0gwhl9VyVKsqAhg7zIUqQMCSko+TNYcDvD
3OadI2EOYNIYD0JIbyMzRDI7wDWmm4IGPuPn8Zyv+0297m3bv2rILuo3oMUqlSh7
wehYb1dlu1Njv9pRcbVKCNNactrEBZWP5gS/YMs0X/1OW5JucFdz0bY4ULFEvgiK
EFLmRNbBDWFluotJ9uQwQU37YOKZi2FU4FYxU4YokYTd1I5g7HsAJRaguA86C5LQ
igM4DImhHtxinuhLBe70WgcfqPj+BIjhYcAfI2CMxKCeIFPkn3i+CcU1quVo7gDv
TrBvc9zrgT7uXpLPvQ6q+0zPjPROUZwqS+GcaAgAt51GfGFoQjJkKc1XVJg54xUh
sQ/NLR7ksxpKDYG5Z1QdZdch4107iwqNbjLzOiSEKRYNbn8fND6ebpZ49OuVa0zk
dCEP0igksl3MedunXLig4WJQM4o+e9HiB26H0Oqoy2tvclF8uI562gxUHvmY8ifN
KSpXjLMHsO8mgFuco6uzwqFKvXTefl8MJ8yqQquPpHmw+oCpG7O3nZtUY5qywDo6
3RGB1jZSmZxrq6Y0ubOlaRHtQyH/JVX9CL8E4Nf2YHTjMTt07qEA0AEY71YSEkIn
H/DF2z53n7eXtpHYEmUh/Yozh2yfE1aj2HJwxnHBmGDp/kpuKgM0mIsRdr7najaf
qIO9U07tiNw3XYuMl5LH5J2cCbKeOVy1/BZwopVUkAJTq7hAccHM1MP2SHr8hVer
mi3Fl21gH5QHfslF42yvLaQveiWW6Se6z+T1DL1/m/bPHiT4lztMSb3ejfqCLvRU
S/rBOV9j/4280KMligosAmUPyHCAY9V/0VEU7PPH8rD3X1BWAk8ryX7BtpRzh96p
/ld2Pa9keAf3H0G1HtqQHRlOTqBEPiP4P4VVe2dEHgHHtS+eOd1OmmYhtRdUta/W
q8Z1M7kVBSEVgd+VOEKPVpIoChoe741py1JR50h/k87xhnwX7TArIGKQq/aYr7Tg
cstuSgiFc3E8nr6AXINqzSuBp2aFRJ1bR7bE1AGmD7lb6i/nbx582x2EGULpeOhy
olp4EyNX9ZlF7xJnmyRHGybnGwZuJ4iQhWWV+GPYXZ2wcwqiZrCfjYEGgru8v0WG
rk7bWBuJTg5RN/baGG5ci/wT923ywfkv2HCbx/T6qJIqr+VdL+gspJz/Q0/zG/Fr
O48TGIQ8HP7pjSuzaB2woUmkCRvck5fJD458HVysy/Ouzj/7Qfw7ycfH9htA9WyQ
KWvUqjwrBiqI3wCbfViDu8V7GBFyiZYOHX4MzRVUUkva4NrycPIu57fPPnPR1FTS
1Gzj7TFzekdPgUUmGI9UyZt75C7XVKuoE3qPC737XlesmGgayDF/kNVOvmj65bHE
vBQqJk35Ex80D1c7ryzT0ehHX+nh8gfidgxlqUcJrOi5Gk2i6zWYvX7znEU7abnT
9Wy7mAOAmKmav/aNVDpVV+1mNq2d+HtEhqulKjePEGCEkG0lF7VCCBNDA4Z6heHC
N1wqcLXj+grvLdTMOlNrk3CdGP6I5ADFD4stH89GnrBS6NzZmqBiWQ2minfdP/ye
+bCEEAUPl0MUWrIYBioDPD1EWk6qH2EeJV3D4jnMehemqJx8xLdVi/mADukVN0cx
P9yoOgb4dQAXf860Q5/dGmYyirGjmiZbW1hgj8lizFeAVKgGSWEJCSqCfQY8GU9f
v8llbWFsQpzKWFc1cByEBEHHTSOZrPKTzvSOk9A7/Z6eqi/n+0Qc+wtPmGEiFteq
D9bO/8W5uK5OSZfTKZ6nuhPbRU7oyEV0N1UodqJaC8ebE+HRFvK+QHzmSZHygKCj
/+tC3w+mJGpc4jKiRfasLDSMlQymf3xLJ60pL0+7bLUJEZpQ1rta/LB3Hx9WoyTa
o1uLv0+RDuCFneeHV0ChIUAJKC7k15DfIg6ei1l2SlqccV/m7dXQ00GwQi0d3s+L
hbARALv/TpSasHKT13pfcZbTCggs4/f5/7c5uUSuY6jvhYEc9XiepcFWhZL2hKgZ
WHNg25tw1Knby+xbdyNk8agZlylS7Dt75lsMS8BY3KqimIWhv/PCsAunT87B7vaJ
rKIZK6kYmy19IGrnW8m2LWDGeDNo0tfwcBEjO8hEhOkRy4E/D04wkSVT4tYLeFDC
vEuf6/4zDTiCWBS0BXgLvHdmJYqa24ZlkOfnYRb2noQ4Bz2okg9daDLtPyukoQRr
OiJjWW+/adK/NQviNVNDlHsNwn/bB5McTD4TjyXSfh99gtccoX93bkeOAPRONfee
tR4TzMCTIEGZf7lci3OlUjAMPqX+aYeM0sUkrkHLTUFbsJi9gOREJESaZ7yjw3+c
DSDxPSRUxk7i1qh8BiK6XdZPKZVsY37I3821VvrBUszCR1chG3k+fJcInyi3qgyY
jeqmMB+DyprLvYpSP+ncHJZxB2yeOSF0kGqUuVScIcB6cpOGwcg1XYo3yrhJnxdO
410PrEj2/Tz+SkXSVHF2sDRF+Vbm1qwJHrDdMvY7G1q4DdFbzzAbGAtAbYoLWBy7
uPJVJFWjmmw5T3FcXKk014ozHe1dem5CG5VqjKmWVf6qhb4PNb9XLjojwyEFslEl
eW9WD51T2ic6CFz2yk/hJj2lHY2hFZZWs/2E2+YL/U7h6laFld0v9qbS07JmNwl6
ysRy8xq25H8LQZpwVd3ru1MLpx7mNQDju10BkT7M2auWwYvzw1CbzEx0I38QEBc9
hKyNpzrJD+PCBkcMMKOqVaDxeQDfE8JFtnMNlMUaG9Qv4tovF819FDPtXDh5nFQe
HjkyKSNlfi35Gp/w0cziRInPTnrup8z+GHrmtP6hndrVnU8vgopAXxcSlyAE9Xal
5RaFs7eRoexVkHOwjzLiknwNlDMvwastvzJclRGLrxG/P/ayvfQkxa+PHn9/Aa1g
mHT6DM41Gz4KEjiCXZfhITwRYJqSR9Azxv5L7HBfz9bhK9/5LA2gvBqB9NhHK3oF
veLYKdxAJtrsKkAlFpkzReKkHNv+DN0b3yHqNiY0YB7Fm9XtlR81wcphDQnwRCPF
IJbiLp/Ft9AMVUfedL1E7GQZiltYdCHDwC4h1+Qd3oTjew5GQt4KgfhC8JSlaQvO
tK9IOlkGTn8FeXtHqZcZvaYwhYRkYXxj2VhXD4L/MkqRRoOnx9JNN0FMHueVapsc
WVpv/uqZLruossarPxnvvMaxRiic2u3jE8SdFxRMMbnjhEdmgHz+l+bGxDMABMsm
0OhOnx4CIHyByFCYS5DQoIk317CYagc7ZpUVe4wN+p27wuY05g86Jd13lDmJTIJ8
y2Rv+VY4TFcXf6sXnaWxvfK7K0JmKulPeRnxFo7Y4XVpUnMW1JLTlDheNjoJt2dI
DIXB6o7390YHlcJYHd8DsMGcxwdtNtHRm0SzNVQ0yt+pRlrrSZL6S/qgv8c8iIbi
SEF8W8g+KXl8T9B7RY64wNIRHTCIcTIbWDbBi9KoiOxPMugSRPLdbzdLuXwGuxQJ
ptE6kqje18N6DF5cn8N1jDVAdQLRpweeZ5QbX6cfZU3z81crQI/bLg6HJIxnEClN
XkZu4nf7RuRCs+R1J+duk81UWijnnLm1F73U48bdRUEqTwYURRCLBGZUp0PRu2wS
1HNTCKXN64OmlrOqsiKU1kollwOADsclj1DJGpFKmVrzi3bPQ00yYHtXH1+Ktpym
UzW9lhAxAL7i0GlB9voNu+a6kGVvm8JyB6KTHSEfouvY+drOl1YkBWmdyWKIgymZ
RaASkQWcFytBsUyfWxqfkLynsqd9wQ7frOyfYZmIiDpMLEJ0cR8jsmXL8P8Q5QQS
ksHV9s2odAdQmLGrefoPT5yQcL1TcM3IHMeeup7PsB9E82ob0TTSLnlNvFQ/3VG+
MPcPLZ3IQ7KaRjqwNY3V35gsQMQ5MoGRklpofHYyeZksbSIlJqLDirfsBNpD0Ukb
FC5kJXfVBBXQ7MY0hjuqYbQS5wcLZxLvcZO8nrQkZ8sgONbWmbx/M9pOdyzYTO6k
YP9oQ6RvmMBU+iq2e6caD7uErbpFMIFkDesuk4iwEYScYlY8nPeQb+D5cpmZiwsk
aR61+FyRuMDODewaiq1AMtZbD8czi+jrc9gLafSmSQWqo4lsRfU+ysbLV5c30/VR
fNFVYubQXY1YGSZb3UT0HjSCAgsr7NbPIZf4+cfOuCv4m/BCIIMSdd92+i8miw+0
XI78Qa3/h4pWA1bzXGFYzHMTy4mFoA2mATWORg3LM+FGrteJd2I1qD/wL7WNsqSb
VILmdWbUMhfOxC408nZbTMH+j2TfCajumGEBbyZyu3zmH4SOaaadYCSA1pxryLKR
O8BdVYG2JNZfpxoWK6AZQYH6sY0vXiNvPZXgPi8ZJmAqqjd7ed7TBEzPpY0O97Kg
SxG0IcY5CLyN78OPe0mYRWC5JHIxMk6+LAuPv2S3AFe6VGvHRocV/OlJGLIh9875
dhr72KClMdrlBjG0mqnsFhRWPDwYDWwYCNeZcRtBixoaSC3WNAEDkHx6M93axH7o
BH78cwZKj82DIfv477FlUpjx2rCfHp+4mhOpNmlmwm8u21sEJvhyM0GXIWuIg1XB
QEv/RmWpIMKFeX/xQEhx8CLln8392Te8DAAiruU+Wide25//c6gNvtCPmrXiDBOS
+39jDpSq6bg76agrAamWWSSYenSdFfooJBnbvywECqxjKZTbmDKGHgfQ0r6mysDm
JsTEMEhiC6YP58x8onvIbJKUc1QzIj27+mvB+ks9Y47dE3RMu2A78Wo+J4MMe1qP
q1aQO5ht67u1idK8MEA/SllX4iMBrW37EU8kKS5uXig4XP5UOM2n7fWvGjivcnkI
EtqLeNAHvCLOVkUkQTxFM7YaEsKs+lDAgkvJM96fP17MwBi7o+alhCnrnEwfUDjM
mZHfIUqMuOE2umnJmwFIrL33PAfvUDfMvC/RKeLFr7MKleMExkqEHHZ0UObt/QsY
ZTytKURwF6yHUmpDB6/7FVRTbFISf2MLRJv87y+vLuvoLATTeg6NvmRjrqF7gEYp
e9Mac1bXni4ZFrKk3fLeL8vti71ruN8bXYKduyvbJvfE52zAsbBFxnDvHbA7JxOs
NA36iXCrPNKzeP5Kjcns3qDcb5amtjcAdr40dKOZs7WmmR3d/l59JfGv5kpGQlQn
iPeZubVuimUyc7kIQ/eiFe6Kp4DC68cEkkzsx5PZDopCE/UIpzjjZyUC0Z1WSU+5
4wt1gCnRdSduuu7IkHqbH0UCc59pxxRLKMAvT1P8/5MW9jy5+mSL6X630qb6sLpi
k9KPowpAz8GxCoFe+UUdb6Uxpk0UacXgH35z1NJyVcyaWrBiN5RGwGOeykwPJe4I
hswftwE1aAogWOIsSNAtOKt4V7nKftOYaymX7GcmfZSsbiaAKOpOJDz2Bbtyc0f0
UXd8pxvpQpXdsmr0c2nutEr6UbBmKwhMTdWuYlOERPAzrkKgXvNGj9viUB1ibwkR
Y+zIIqvrhcC7itVIMXEqXbXu1nh+RFcnVJ5y6XMpIqh5QT+A8KUief6mMAvrkFaZ
UzYX0XoUf6STXJ1+pxHLntF4raN0872dnN6tkeDMFUxoDDTLIYkMYuzgV6EVhH6h
WzMwU0dnUABgng71uxfGTxebpQ5DNKNBt8y+vP9E/mB+483WVWGY/SkCuYLcijVX
7F18+PTYlynb+ZWG2wtAEpq83tN/Lbxf36r2aY64LHeXzXsMmW/lyO1+GQXLXlzN
icMUP1HgpwTFQ7XBTN0Y7KFpP3akg6MiJvuUaeFktkC6KJAK6BJSQ0q4bIcCVMaR
GWYI7dY8ybsoMPHNv/PuDYLdwrHmJmVFO5YT89slKScmkUpTyc4YDQO4WsuJ9cdc
EJ9Y+vpGy+X8y4PL0uZx6H18RONWEKeANxtJWHPP35S9hB8WNzy7Xo9K7YB5830H
NCfpenIlsYkGjg/zZ3IPrZBWDM9m78zEPm5zMlnSyIi3gievSjfE91kjFWv71TV7
pLuNs+bqnAfUqQPiY59GdywECk9YLIENCwS3VNRWpOjYHMpEeUTSZIL8AKVCRJrM
+3MDgKhvc8ljIeWvU7kYZRKBKQSqlNeR3TFTmELCY0rP8L+ruk1NetcF5m/bcL2Y
EajMpWMJuVOD3aIOT/qQ6ez7OuC+8k30Uir41DmLvtxuMQkgKLPFMwB3vODah8X9
btr9QfzBF2emg3XQqOlkGAwA4Hcuf2RgozBzFgMPhPGaNHZCCN77cHgPd+EajVNm
QaSkrF8D/US21S1HxEMsnVOemLgzmcOyud2m6AAv/X/hoeYUHOWowG1HnBSFKsBS
tSalalVrQnSY/fKC3LPoAdPdwzAoSS1Q/fWlTjgGZKeXalhZWPTVYsCqKMMzLiU9
zZrtvNcz2xWKUFiMX2/lNG9GmMg2pB6oo06OrQ/CD8Y/VMxBD+QbmtjGjUcadlTO
TaYf+CNOvk/LKbbwDfWYculTA/YhZIW8F8xSYJNrDW+aMOiTMBvMkKGuy0Tz+j9t
g49uaWIN8YURDHqUYP5quH7m3VUbPUCkh02e5iykpIyK4aLntgAMlwalKqcZkhdw
NeaPJeLC8MBe+C6SviT3svmVsEqRrMuEw8bjMu6t61Y7W8bq4b45QvPBER1PdFOR
xpOSkQkrX0MSwTXQxTNjxIjdaw3Sx//dFw8jQhC27z5BnSK+4RO1HaAyoHI/CEZV
98H/Q3U+SEXEfqj0J4ogcxYgbiXjpTpp6AtCTkSbXv6WSobz9w0kND3abt7DR8o+
hNzxfIdCwdjAe9TR6HsG4yLXV+uvRPd2Z+ELkBRcmcSWrUXbVswVyb1oxbLvGhOR
hfF2E5Kbn8zArm/xqoDu7UEoCOwUwFRaZ9zAyUU+fY3XFh5ISxwoe74inrPKv6hS
R8EFsqaP1yTNmDhX6whawt/zNXv1eK7aSa/trPzwVrEs+kgUlSWjImQiBj6u1Dgr
sYxpAamJHcJSTjoMY6uhHAQ/9InqYegKlLHKdrtQ8n01pyeeWtCjyq0QG2mCc3Yt
NZOtDIaeNjJys2Kv/HcoedqkxTxoRxjnPNrLpPA7v1dHVgjDhiROc/8eFGL55bt4
6xrUU+FcGYGbe2Q0thakjv4pcktEXpD3Oing6eYqewrFmB9eWXUxAOljfvormFz3
Flvv2EJwIxymGE620TYfNmhZ0brUsxz31vI3TXPJjFwj8XU4oyfKwKlTzTnTZMgQ
fITPijPK/LDoQmNH57vUnxAZLYcOvZHOOvx4vlzfK89sfhEt59p6pjv5xtMEJwWS
OMGe3wsLSfwYnanD6h1VpM09L37s4TWEY+lfv5V/NL284akwO30hwuwQAqfB/Aqd
ViHfmJl+E/NXxwWJ2s/lchD+H538mpVAabJPyh4JgMDday28ksstAB/oGLEcVp89
rnClAWmEXxqDuiHqamsq7xgenU5Z/IydYSwXFknw7vG9iQHw9AmkGXw871h4eTTG
UXKFE3JZLQk4WLXaBX3qBSwfBZgfLayJoBBcPIQdg0WgUfK+P79eFYguPA3XbXW/
YAAWN2PESqot8L3IHZbz8WLR+JrRRC8WlAsXgB5aLJ1eYMw2fwvNCSIiDiJaacVt
XAHP+427OTw3ZQX0H8PjBNzwKChJpGwRPXi9qHscWLWKw1dhfCLGXy7HZL6lWGPO
50XPBGoOkoiLC5BxvSxshYFh8peZ+SFYI35ejLnQtkBNFr2OiAFYKDEYb01Zm3+6
DpKr2c6fVcSXclo+vaIVeTc5TB/LIdZn5sa4spH92/pkIt8v8ZC22aS9YODehURu
0jcl4ap7eN9Xc5zTFktUUHXEDa6dFc7mWscdJt1iMOMrAcSXt1slRgshbJlkwBVz
p9hNHeuBrIkUxkMVU/YbQ5yDztYEaBYOh8HIxNgAkUFf9hT+Gu6Er8nID4k4Gmk5
BezrVSTR0k7pey4479Hkm5dqrXmEIwJGv65+BUvTaEj4F+VS0DsRKAZeMDdZzrAY
hV0svtdAwb5EcI9sMgDV0ETTj9tht6eLAUPU/TZI67aezqlP+1pq7ulOis51j9zE
x4X2ajgQ2MhXBkWV4tuAPv04B79db4M8LcexnUZk058lhcnmEwokDvggzJdbJo99
RupUQU+Rt1+T+nY68wEJxWn40VTrp3Q4c4xAN0d/s9lECuBpb+PLassR0iYoXmhp
Zucgs0ZAKs0+BQpZq2Y2lfU7bVg6kOoSWrVmLIRwa4IKIWFoeiTGcLGDbiYmJMVz
zfyIEqxSESrNHA6VHXDc5xj2gxkNNPr0r6d/motR6uKNOvq+yqQaHOwGoQC/K6y/
fitEJsdKIeffuAOz/sVdI2YnXIEtbIUOVcA60kcl1CD8pgb8D0rBrJGs27f2hGoT
eNtND9VV0MZ4ehlJ23gX/NIcdYq4Ga6dY4CjQzwsTY3ay5PnjlbaPiXBESCZ0Vr0
5wYWsshzuA6oobilVrLwrkp5kTIdgr/ROkjIO2vstlSevfiSlWkXxiGOhjgfoXa3
eiK4VCwiW7WdYOFz/DzK7MrYCTn5kKL9kDz0TvdQCyR7+tdZc4ln+fKP6pWHvQcm
7uS3OhpF97mtQQhWS8tRVFSeklrmLiklm+2Xry+pbthZFND+oDRNw306ahhQWl7B
uV751ws8OzdJOtQAY/HlKkTuDVM0Lo3dFIKbSTe/Q8KcVFF4qbOb87IEMFpwQob7
4YeTGJBST6rz5Xu3fsvljfLZB6+gmg9IeKFJIDPwmK0bEVPh6JFdmQEYV2ChDEZn
vdxsiX83Qmy1zq4tjJkxmX8VPom9Fi3Gl/LjFuYDzKr/jLnIXY5hDZn8CNzpUwIY
6SGflaU2CE3t2WefzgbZm11aYo2bCRdo+2DcEAG1YKbKs7dVUJkvXqGGGeViNN1u
W+x6Be5g669XbKG+Fk+RIaMPukthiw7SLs25zOv9w0bZE62g9w2RIHLvWyJUzJDg
iicUDiH/fWDVj5CZDQN0Hiux4574lY3fH3GFY61iOIJlGflex5rTF3Nc99rqYwST
MfxkQmq+hrFn0/fHideMyxQS45WVFFbpQ/VKrwYXDvcfTN3V1E8x8JvTnInC2jUr
164pvHGBTmYcf4OwqB1aPVTqMSMlR5EejQxFMxDARYOG1DwWi3b8m+TdbGyod00D
dyR0aSyfGVBoygXap4Bt4O+d2atjMcnB/vxoStZZlVSLckdrSBGthUjBmnehv6kN
h1Iw63h9PlGJhnvlx23+9HBR4jSb0+vSZhph6wR5WGV5kRAkVCql5CUKue4dNRv4
lxkMRHuPuFNvml164Dg5R8iTDyqVAzMbAyMYzUI7tLR/BdL5D2Mxf6IlVUrrlB/V
Yp+e2AF5xEUcYKcMSqj71RT+hsjHGcuL6QULk4OoTZNsQ2J2AnpFqshYeAfqSC1S
YmlSA3dRh2OUxe2O3YZM411YPNKYeUqp0dPn8MeENaeVySV2GkUkRKz06f67WcLz
s++XfWX6rYln9RCHfsvo57mv+AjlEL8kGuZd3Ueol6RbLndVLx44r4ZVT43C3WkL
boc2b4D3UZ8a0VKmeBie/zrJ6dv/QHUyWwxSOEgGwFt3K4YIl6zcleewqUEWRnAT
suNbj045Kpf6e2zOnh17vtC38ZPnZVgdPTRxYvIkE8rrXY84Mh9MUHJOXCs4larf
EIdjwEWMrab+Vivt9SYpcFYy7sGGtAqEg+c+VfQ+nwkEqnx9vo9YBSYRoY1cZcud
Kf0EAX3xK64ga2u6nSD7JKAJI0Yhx/BJRsivxMjnz5Q38Qtx5PrLk67RqIj+Qgd1
bzUEvZCD2KqreGravNn7DoTwDMdaqx3uNTg3zzHOIFhpmOwBBHadAqkEJxv9MKk/
lCYh2Hl1b0KlFPfq2JibbaLDtpa2yKpYrqlyBDX3EpLV797zn5VtMp0doxA2ZxfI
rynM39Rfy1YwNBwnivJTsNcw5R5ZRjdCar48MqENwBy3KK6zSnoyKbdktDtr+0zp
RRrRIQkYhxDqhDtzrDfFDBI/+L81UvOy51svGOpvAmiERYDeRgKO6lK9I7kIOqsY
UKX5RTvZmhaMCExvK8pcEUULxM3DeTHBBW9xxvY/6lpeJSryDL5mslU/4A7pNmct
clbTVexbveEPlsHdx0c+GyDYascpv9KmA4S0rwrpYw1iprZ+0q+Q/yEgz/x59L/K
Lg4ZFnQWiWKGj1QsB6Nke+W9R7EoQyKj502kuKl8uPC02wL35R+8RSN4fJcuSwuB
IlX4ihhwrdDqW4KajcLyKW+Wf0YJQTNa8zJpaG3S8aejSc9IPk8jxhCMSPC8houy
IR7FGybDUoric1ocpkiWE45qxrIFnIOID7Um8q2QOvNbghi8Ikddq1xT1kwK9l6E
H/A8Xcd4T70cCunsRdu8vJYvpAmlSEonlTuUGCBN280Su9oN3tELmae+/aLT3rP6
Y4XTYZYDStGguoquH5G+kTqc/SHDQCmiluKtIw2/5yVlmvx5KLrGtaXwfVQivxA3
tL4jCkudIh9EKPyReP4pYUqrq836SWGYqL4Un6i0W+opY0NDJRQnMtWtAPiV7+Gm
9qZtAiOBB2SiiEz8m107WooP77fZYc0zsGo/PyMU0v7ltwyA6/gx5r8AsC5QxQQn
oKBET5smim8K1htBmKk72Jqnj4PvrkWznBatEz20nAG7+HWpWi7vovS10sXNFcgs
yi0AYIOySUGKhDdv8diDSTlBBioG74S2tRcfqyW8WEiwTMf411XP/PhRScEsrsIi
tbpRAvh6CjyGlU+Fm5Q1vXBsfvfLiLFF0lHH9lJJWW4ZzRu9TWqMXGlcDR6MhBxB
KcFTBmvu/utFOfAYpVgO6CWKdxh24H/WcqP23yDVN/+bkzG67a4SG1jfZSsTYJ2u
Uwf7ACh8A133i4Z6+gyhtQEZSp69i5fcG0RbPSfV9yTiB/LKnsGqfmCbnESZNnrq
ymmI+OWJx1WLKtuGFMsh7apalqw1/KScHoSX8VGEPGQAn4Uz0D6bIUxOhgUe9kVy
oJyD0BotLaPPHSXuf6O8WojYYAMS3fgB9OIJ12UVWblVg6JCrwg5ToRDOlT1yhMl
uqsCCaVpQWal+0AjEB37vHPUxAvuHAWOg0/GxNMTRp0brrt2FFShp0N/3EfUptrK
L1O8IBSy8AIKeKl6HT32QViXu+6I/Ns/NyzhNYrciL1TDOjoBWNtRkpZqGkAn6L4
mK9XCza5vaNDfKLNtCOuLq6N8pBrFbUQdZEf/0VsBe7H2w0daVkfMYWKbPOq6QyN
kVMr4BApGirJj7dYMwka3in0b68VRo9rZPW1apgfy764DaYdfsjuyC0s5K64DBOm
nDMSlJqtnbfaYBl/pTQdEZ6IjKO7eMYVQvP08OLSihKdr/1lDmA3nx/M328faHdE
VFrnWSi/AfZtqIXHcJyN7o0+t6hGXJacVmMFhkvfsmsPtmY48puDL5N3lh/oJfeT
YrmBysyhfQuzKQTiBNdYxMzr3fF8ebhYI9n6vU/nsSackwEmg7fGADWA5YfMEm2f
cuRK5qmA29vV4aBydpu2v2b6XXSQ5iw7ElWzsP9aAx7z11Vm0z79z0rvboOYu6LR
YRhXk5WSHxrxEdRtjB4hVoEq1AMIqPq61VW2A3mslR5KDKMMR84xy90iciCISoQR
V9wjK5THwEcSpUpuaNMBK4nOu7FWfiyGEfciYi5CnVyr9VdPHb4zA79Qh3be3zaf
ofT4n5yDfxZaTCEkjllXnyMd0HvmpJLOSb/waI4gskrtnIwMdUp4YXoezZHvlyvs
T2vphxhvRjlKS2Gj6s7HXRM1jJWRuKf5v5N9ppfQiEQ8JkiYZIz29OgBAPj0C0f3
ZD5tNhxfNta01dCb8//wVO+k/oGgDTUrNyZrS6L/c6DupvwaAOM7pXfXojgyn9+s
hepwg82n8fXk2SLU8CiNCRXGupfaPBXWQ50PF9c83ZJe2eYL7GEPYS9JA0/jedGv
zbl/U5l5cbt/degWt4ERB9Jk5hSSZ52WdFxj0KLFePBsJWj5POAwioKVQDYsJLAt
qWr1mo9bhc7BvolznFKV704cM+ErN1IhTGhICwWBVj52TNQcTq269Y1FJKCQFRhC
F/nJVN8brHk/OJHIaCetgPSTIgacnEOgzEwIzVLYgvp7SiqNC62T0sK9FelD9lZv
YdHkJK8YONYZfvedyVIuuDquFEPjAJt71bjpUtMHJAWGPRy/VxKe+ryeOIH4KppS
cB0pRK5AsmtTFZMNosyVpOUDLAlM08zEQZg+xLzlpFkBFz3uutZGMJVjgc5vW/2x
gVbdUBncKEsDLiwzUun4tt+lpU1eIB/QaZjDMCUWLu4=
`pragma protect end_protected
