module q_block(
					input        Clk,                // 50 MHz clock
                            Reset,              // Active-high reset signal
                            frame_clk,          // The clock indicating a new frame (~60Hz)
               input [9:0]  DrawX, DrawY,       // Current pixel coordinates
					input [2:0]  roomNum,				// game's roomNum
					input	[2:0]	 myRoomNum,				// block's roomNum
					input [9:0]  posX, posY,	      // location of qblock - will never change - ORIGIN BASED POSITION COORDINATES!!!
					input [9:0]	 mario_x, mario_y,		// mario's coordinates for collision with qblock
					input [9:0]	 mario_size_y,		 // mario's y size for collisions
					input [1:0]	 is_alive_mario,		// is mario alive? - if mario bumps a qblock while dead nothing should happen
               output logic is_q_block,          // Whether current pixel belongs to qblock or background
					output logic blink_num,	   		// animation for qblock blinking
					output logic is_empty_q,				// is qblock empty? - used for animation and for qblock logic
					output logic [8:0] q_block_address  // outputs qblock's address for sprite drawing
				 );
				 
	parameter [9:0] Q_block_Size_X = 10'd159;	  // Qblock x size
	parameter [9:0] Q_block_Size_Y = 10'd27;	  // Qblock y size
	parameter [9:0] wall_dim = 10'd160;
	
	// States
	logic [9:0] Q_block_X_Pos, Q_block_Y_Pos;
	
	// Next States
	logic	blink_num_in, is_empty_q_in;
	logic [9:0] Q_block_X_Pos_in, Q_block_Y_Pos_in;
	
	// Misc.
	logic [9:0] Clk_counter;
	
	//////// Do not modify the always_ff blocks. ////////
   // Detect rising edge of frame_clk
   logic frame_clk_delayed, frame_clk_rising_edge;
   always_ff @ (posedge Clk) begin
      frame_clk_delayed <= frame_clk;
		frame_clk_rising_edge <= (frame_clk == 1'b1) && (frame_clk_delayed == 1'b0);
   end
	 
    // Update registers
   always_ff @ (posedge Clk)
   begin
		if (Reset) // move qblock to storage place
      begin
			Q_block_X_Pos <= 10'd800;
			Q_block_Y_Pos <= 10'd0;
			blink_num <= 1'b1;
			is_empty_q <= 1'b0;
			Clk_counter <= 10'd0;
		end
		else if (roomNum == myRoomNum) // move qblock to the right position and carry on as a qblock must
		begin
			Q_block_X_Pos <= posX;
         Q_block_Y_Pos <= posY;
			blink_num <= blink_num_in;
			is_empty_q <= is_empty_q_in;
			if (Clk_counter > 1000)
				Clk_counter <= 0;
			else
			begin
				if (frame_clk_rising_edge)
					Clk_counter++;
			end
		end
      else									// move qblock back to storage place
      begin
			Q_block_X_Pos <= 10'd800;
         Q_block_Y_Pos <= 10'd0;
			blink_num <= blink_num_in;
			is_empty_q <= is_empty_q_in;
			Clk_counter <= 0;
		end
	end
   //////// Do not modify the always_ff blocks. ////////
	
	// You need to modify always_comb block.
   always_comb
   begin
		// By default, position unchanged and velocity at 0
      Q_block_X_Pos_in = Q_block_X_Pos;
      Q_block_Y_Pos_in = Q_block_Y_Pos;
		blink_num_in = blink_num;
		is_empty_q_in = is_empty_q;
		
		// Update position and motion only at rising edge of frame clock
      if (frame_clk_rising_edge)
      begin
			Q_block_X_Pos_in = Q_block_X_Pos;
			Q_block_Y_Pos_in = Q_block_Y_Pos;
			blink_num_in = blink_num;
			is_empty_q_in = is_empty_q;
			
			if (is_empty_q == 1'b0)
			begin
				if (Clk_counter % 10 == 0)
				begin
					if (blink_num == 1'b1)
						blink_num_in = 1'b0;
					else
						blink_num_in = 1'b1;
				end
					
				if ( ((mario_x + 7 >= Q_block_X_Pos && mario_x + 7 <= Q_block_X_Pos + Q_block_Size_X) || (mario_x - 7 >= Q_block_X_Pos && mario_x - 7 <= Q_block_X_Pos + Q_block_Size_X)) 
						&&
					  ((mario_y - mario_size_y <= Q_block_Y_Pos + Q_block_Size_Y + 1) && (mario_y - mario_size_y > Q_block_Y_Pos + 9))
					   &&
						is_alive_mario != 2'd0
					)
					begin
						is_empty_q_in = 1'b1;
					end
			end
		end
	end
	
   // Compute whether the pixel corresponds to Qblock or background
   /* Since the multiplicants are required to be signed, we have to first cast them
      from logic to int (signed by default) before they are multiplied. */	
   always_comb begin
		if (DrawX >= Q_block_X_Pos && DrawY >= Q_block_Y_Pos && DrawX <= (Q_block_X_Pos + Q_block_Size_X) && DrawY <= (Q_block_Y_Pos + Q_block_Size_Y))
			is_q_block = 1'b1;
		else
			is_q_block = 1'b0;
		if (is_q_block == 1'b1)
		begin
			q_block_address = (DrawX % wall_dim) + (DrawY % 28) * wall_dim;
		end
		else
			q_block_address = 9'b0; // don't care
	end
	
endmodule
