// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:32:02 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NDf4qEU88AlXWwPmt6+cKrduqg9dBsMJGlo9+z+rrl4VEPzHkb9eIFoFWox6+/mg
tWtpfZwjpQw4ob2uMaQG58PYVHf60igwq8IeqGYcaI/zoYf1kD2FwrLM684sg4h7
Pccwp2zzR91eKzMoV2KLfjgkLXTk4O0yatnYnu/TYfI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12240)
LD0YYakR0ltLdOONNHg4nWz4NNkFc0ejk8QZabquCjjRyd0DFgbuhkMxNaix23Q1
DacCmLX2uaukh/6TzsFDt3C7TI1nT3+xnUNWchJHP6ZqpUgeyIwNiqusgVWHBr4H
tGrAJTCAgkQ3Dd0mjMUsA7WUqIO1oB5VrTk7z/TAKTQ7aSG2h/yPvSWbxV72uZdV
8OoSnrl7iDUGjWauzaltSLittGwwjPpQmXREjXM305kVh+/PCX/Ix8mgzhZTyY76
FdyNxJyN/QPgPK6E3AXh8xya7GuFZR3m95/Nv8ZxQ8kAachXSfBnTb69ruHLCm5R
YTt+Y1/YDepTHeJuK8SgBYTh0v/IzUqktQV2rli5/HyYMhuyEF/VNcM8NlicMAl1
38MTc7gYkNai5Kc3O3DlKSFxU2k+R7J+xeohNOlVAvg3yk0f6b5ymndjMKSjltbo
2YKgKCRO3Kq8exEuriwM4PXTx4RW4hmHbFavgbKVguvZHrJT1tNkbHq3J5fAeROu
e/okIg7o5B0x2+IywSALBUzCH6qL+MwvSR17jTUvBglwAk/LoAdKAWhWYPQqqiG6
UaUz+jvZ1n/rzZ2Mn6EKuG+edKWLTqubltRKcKHTNEXLgAK/8RNO55myFXsTPkGz
9a3KqouauEkzwK2Xnm695+puKJETtFpbKrQ68IXQ7/YNkcFCG/L8GqK+r5OksSa7
5/WuXXiWlN91VgMNkeUPxTlrGA7+vP1juV04IT6A0grBQRLJmfmr0/hcuPVtIzOp
pDLnUolEK//aIdSCEY0eqewBhwzNKF8FF78bowh2V+yHgK3n8akHQmPJOE+YkhoF
xjRAX/mQU7YI+mhythfVVsil8Ypt/MvfGOp0+Pjm9P3vJiOF2I1L8q02EmakImK/
JT/1WXVw6+OkopfJl7++0lv50REcbZFb7tVyTo+ClOOZN3F7sUIiLf5l9OoDzH4y
xJE8PyLA77tApxbSauJ6plL8r02BfdfStMrHUykSP4k89ifgk2QXKzepyP17CFeg
ytgesl/Wj8SsARi6Jffn++VnZhCy+i4nx/nML+cr4+Zv1a47W0/CqRhcEtKF7Qiq
N3agGFonRJZ1lvmDtkQ4MEFGe2asGg25KYLmfipXCapY5KOi0iImalz3xwkTsv8M
/Aj+FX/pofLx+jrsEKvksMKV4gSOCKRaQVeg/1inlRaHAAHSrAOzByni76AHsMvX
pm5zegZbe22w4UpghKclvE1q8yFHYYc73FVvfsKvl6jZwPk5Z1rJrLRdolMR5c/w
yFNq/qQ5syzUMOkFmiavBNyCepKhcNnWZLtIzQXs87eYFYKoxV7F46wZUtpVLfoR
pgCgdnO2w0bzPKTWs1VU/B89TJN2JXl4eeP/OMereUDd1ZphB66FASBsV+fLIv+X
Id4P1w6je/WvJKiCu7ZKJ9+oWNEND58Ftj34A7+SlLWYRzmm77caE5K04t0a20RD
v/qp1IGDjOu7ThWJjNGOCTKoyPA/y4hVTf8n7+BFqIlsIaPuMZlEs+S8QIzTnwJO
YHQtp2wVDUpAJoqszvBCGuf44pRQeSZe5s+0hMTffMLA3Eky6sLQ8aJpC1FxSCPz
FS5IZvsApAd+yEYhG/KWJNGNtL8VX3YJKsZM683PVCQ7ohrPHBkkaBet8UcuLjRX
QG1OHhNKy+dXYsECC6kk9RGnYaappT2NjF45cwUs6FyIW/f8T3RFQnnn8BkE71kA
hOIGq/ku/B88PUUH1U2REW9DSPpje/kLy4QzYlX6gjXi/TAA9CfT4V+xEsxO9SI5
vTXocQWa/oejUH6c8KPGdDR8j3IwLAVBFljp6VW0XQit2C/OXkJ6PDESz+PS82fD
p2y9V4SfP857Lc/W0nZYit1zRZ/7HlV12Nl0RC/9anuVfTCGo2TY8XgsxUZk5JtW
ZeFmaTwWcR/fJmvlRCHUHIz0LQEaOuyqHarul9Lrvrnar+Bf+Rz4tkLnQdRMNHil
O5eFDq4E8nNcNADsA+Zq2myN/AWvxvPWOZX1IKG2rS65u1Dto8ahU9W63chGN98M
Cgtlks7Ix2ZSDAhIM5pE6HwFRS9U0lOBQEGPFT5uxS2R7CdkYywbpSGinjT1VvZf
9Dpb+Yj59AFmHwfxp7eiqotXWfW5Pdh/5Pr24JDFqpmtP6k9s3R/BZFTcf2yq7XJ
d1CdSEtCosAKj81lIT4seWPdoZI0AZH8wolIQ9UI5WLRgJ6AL2AffHls+2WjwLdq
mBqUWJkxVoycpMfGVgYoN6YJSx7oZJtqr62nMaFOYvE4iwhEFlf8wF9fioK3YZvG
62lpQ6FgvtPx372RJgy3x6pGpV3FcSOOVCrNHaSgjyyoBncLSPtK2n5ZDbOr9ywh
qlpCf+dmxAhppqEy2SeUafx7Ox8rVOZHZriOrq0j5PoKVlYLdOsm8oE+w9l/Eb7L
auseVmrV/Qd9LFNVEtB2Yi7cTvnl29arvebEOAoN2TjL1GZwi+JzcksT5gSqllng
OEbhCB4LhgjoLWdthItBayNJSeKbBJEtWzIjpFYtywSsC2yDF/dAUR9jWySBtX7p
AdqZDwjBLJQIoCLkwSkUOEgRJCSNWNteo7Ju9HfawlMbI51G1ZvBvZsjjutKFMP4
pMll/DvAA9EkYYt1D2vD00iBiqt7o41G0XnYAduiQlMMImdLBsuIKQRu9GSkyY3i
gzqk/2jwjutJbx4mJ9p4PtnMY4pOev3YFCgFXI2UqDT/7mrFOJds8f/Zk6jYzarG
qZ3XvrZHYXKktDAp5wq7GZ5jfT+gXkQUXOKB+Pkx0B/10fTJ9Q4xA8lD3i64ttc2
7yzwwtR4rW2g4MeXAvSZAQxPH/YHOz8+hwUP/NodvQDWgn6IDL5BDCfgV8uXejaw
c48npafjm8gu+Oh6kzDphnUrT3h8TZmc6suEI+Eeo502XI1cDPydPPuj4CIH0kA9
dqgUNtLDm+MFYrorKqRGcnQtBRa6r5S1a7NvMbLlwSMqk6gmuxTq1MbR0AL1ldag
4o8TGC2w6rak0ZWLbjs/7mi1zGLJZBI9scFBYGBI6wu7QEKULhCPkSuLAsoOl/8W
fBXws4cFKE9Zu71PoG7WDUrcY9H2XNbJNiVrNcghMymQsUmgquBIofap28L/JFr7
UGwz+Wfcr/awaKsfPnmJ3tUATdbz7DTnATSIz99BTwXptZ3jv9UBBJqpV3Z7lJ/c
imeTPtDeFftiu3ZPtT0pjxUY+8HvweJb2LkiYtYgAHvJAnP3R+MQZKBrEim7pqRF
9l69EMx+nh7Bw+ezMtcToqaWxn7Nq9kRrDvYv5ZiN+jENdV9jjuSBBUmHdWBs9EZ
HUaOwqOwv81rBNTo5JMvVUJJIXTv5wwgOzlUnF2MPRN0XvaV8OctijKB7MyPyb3M
Y02+g8/6Zq429tWxsl3Ha3VNG5ITiHBhyCerXKr04Z9toU9BPsfZlguEUZ8QhGRC
8OL+AyTdOIo3kBhlocZr+ABxqmgBUrMKe1gSFnXF1V9zfqCTKokb+nQ5Ub2CPNUo
zYHhAD3H8vC+nqEzKK+SaaspzamRkCvC5Hz9wOsIaE5RNxykhQXC/g2Lwhb+Dflw
9AORmfWYbEjGfevh6yR3U/aqmlBa4IZukzvVbs8jSUPNfQFRcp0V/V7MlfSe8ptq
HSXclNRIVhutJLmQVhX7g5LfE0IThM0X3ermkiENCo1+RdqOqkOlWJYCQPvR19OE
6N66Xm1Z2gej/lTVJOO6Okc1Q9xq1RL+0qPcYzEmtwYBZ8rQQdm1KSFszHA+koYI
ZBOkosANRGrYz3Ryj5gr0PAUlcLUpBpSU9Rp2vom8Els4PKfMM5DLxXbA2DM5TDk
34bDInyoTM3a78yZt6KsRjcSu7LlbiC9JIx8Oz4SOKd9wB1p7rKlzJFFqkctBpY7
x5GCx4YGHRekuarpQbywCwbiTkdEjPp0qBORqvhdN+yBIZM9jw9VXrmrA5lyZL96
8djwDSNUjtKdW4XxlWdtS3Kpi90hPAMhBH6Qebsf50GhxEec3Gx5/8M5JSGqRPZW
ZYW1FKstC1OPqHMBUMvfJBdBX3y2yMLth1ueBJsatZmMHchDmPpftNMNHXux4C7N
84hd47FSL6sEYSEGurHOKcTlnua5FmeU8d6AforSAUx77Uhkd8i7JEg6HodRa9T5
jEzP2wAMnAJHgB3gO3PTsd2vopk9tncXxi6KowAZFasXxbvx2yIZoHJqctyC1CiG
r2HYJ8zZXYMfd66PWsyg0d+dBjpkqHIbzQWVbc5bcbrFHeXI1oDLDNXXpshX2pZJ
C5mzINtE4FeH2P+CHVK65IzB4Q69KIU0ZfX8O+oPLzo/w/ECd23OtbRCoDZfpxfg
M60Tm0uCd7kuPkpVz7HPh6w9vLuclow4Z+A73nRUxJwZ7Ye+c4s6Dhi7Gp0iLo1q
5X/85cLDwWDY1A5ygjClq8D5PsJMXaJRM4aZWSRUlIbg9p3tnojpOW32U9Y0rEeY
jOyRVX2+F3fME0TWL2B5p9SYls8h4d5SAcC5VFva4+7J2eGvlhof9lIiSGGoW6XN
T5rwAfldQb78r0HRukfGIM6O29Z63tFriYCJLTdSoQVsQ+ihDTTpSoi8Lwr6t920
W/yHUej7DLnS/rraKfTUEY2PY2Q0z1UnC8VBzfUi2B/2qOQ94o+7X6Wi8wHclupF
qMg6D6Muo5UPB+piAUb2OXW9ZDPAlv9pdO1qOHoEhP1er7glLA7SlLGc/RPR3e+h
4m79RFVlNNmpziq4arAKqRRtJfQkaHKGN/Fu2sBTxDGJKRDHLq+WPTdk/rN+Bb4W
3TAb4ZxsC60ggISy1E+EgUzyK4eugTptcZrqfDtGOQVfWIoHKbNA30Dp/25kGIWj
SMmZCEkgWIXOjFn34H9+nM5mWYmqVdTATy+qpsihBWwVFISTkCbHzLc+pPjIES0W
Y7giBASNjh77jIXbSxlQWytApX+X9alohD04PfH2iu2kZcSkMV+zHriUfnTl9cs2
lukf2EMLcEPdrsp7QpauogWujkRVQbZfKiubAVqrALgLRtDqF2Vphomjs2LXtCMm
52gLeHaevXPzvJPpqLEY/rpc9hiPfT2vu6m6rJ3Ln9V+RlCiEspw0oOMYF5+aZEi
LTqNxhMo3qt3wpgC96NVsEskpo4SNf5rLP4dlR2KHCgem0pOtU40LCAz/1OeIKEi
k931r0Kpayxk5wL8IrHOzC+2ge0cD5ZRmgkueRGjlN/vTksLwI5Ct25CHO9RMQEO
FrNkSCwaRI6Vwu/hptiYZ93SDuoffygNM0q+RQd4vwVbkJmvOE87L3CHDA88GdtB
K589g0JauOd8h7i+7i2EUtVNznX0FH2aSNzu3hYa4xxI1R3+Gzbbvyt7Sb5Mag/H
mb5wqoYBu3+HTgeiFkSi8fRDfMd28dcrgrXid8CTngWoHVWyhlYt7ywh+Y0GYc4X
yCYbfmuR4UwqjuOH2ytI8j+FghQApJasvkfn/amCJItldMY1UwvmI0daYlDgMo6F
hdHmNkcuATK4Or7GhAM8uwmCACkQ093CUZaQVMqqCvKot9OY80sC4c38bd6jgLWA
2p6igz5ZOlSBgO+Z9iWHZKMxiR1N/tbzvHUQUdBK+DWeXiB9E8PR9fJB6JRqhV/2
fCKsXVgkby2dt9kd/03NKYBvXX11VwIw8pyCIhoY/WONDr5swjjq1SbJ5afk5mg2
vB+G3YLtxrmPToEGeYnMoQrej5hubsYbJLyGPkG3wUA72k/H3RXk217CYWtc819S
LQL651f1wH5q/d0dOMW9nTDKgmKUbsgWeIoYxs8g/xBsM0tfJayI0OjF0aw/Q2Vb
1iEcoD7LK/LYcUCJe/9xzFLywkZ6OsHWgh5EPPhbzsQR03aZmRXMRtiMWcn7BjPv
C4YqV7YgPnT5SckEqIl1ncdTyDsFMmffmEfDVz5mbc+9dY1Qy7OraSkkuhC5cbCt
FL59IxAS15xZL6nhoHjKLgHmoe0G1X0VWVRz+bSXIqarDslG2ZskMu6/2zQ8QH5z
7q2fIVHEeJePEFATvRTK6BV+HCkMIQue/MIBuKP1eeu6xhvODfHI79uHzaBfIUT7
xQQEutZR5tC20n8PIrhaI5jDHNxYHD8wgZYmH7Iu1FYG3pOU0LHXS2NXrJPvg3Dv
s2JB6f2cQZmSCo9/PwrcLtEhUcjC4ElD8cVunx9E4GDpLx1CwB7BaESS4u0o+1Rr
jJ8j/dmXEnZjWalz2Xhb4xdxlQab5yjtoboeRbp3kr1eiJkBI6r7wEvgj3Kebqal
K7MLb/vNWCkcqjjJlw8sYSc5hUwvOwAWqPiNYAMtzHBUfK90eMPcO6rCxbhPsZgz
CXJWzLlLxc/BMScN48WnaqDUTz6pyVtGvHXPJPE0EI++l/OiNzq31d6jKXTJZJhL
4kAlIgqwSh1UzIAEZq060fbMgnHqyng/JuyeEabRj9+MoAqM9XBKhwzwqHviVnHy
1n3nRfCb91Yx3g5UEA/RgJQzFiAfQVfcGqGxO8OJNZ/b4SRWQau/A2JVsb8BSGjB
/nX8PVjpvIBgtDjL+yOIxjQmpM1ROUF+iXnq+EJkelSQibooWZ2W1sGcttTqYdI9
BzGgNoc2Hzqjh6A16pLpYmJRwsNg8TT/pb7X3yxHE2pSr61JcXrfgg0Ui2hE5sNp
EbSThHdyZ/kkCyrfkCxKEmfDFDHbmmNqut4rlNZ+TVkIu3riXJtloDpc+9QZwFLn
kdcornlKI4z4ZFW9wiM8okJYEQ+FhfNIzXiFJ54Ou0Jg8MnT/Hl/tgWWJxf0Skss
tNjShiumfkdKRpBbMZYFsN3OcAtmd/t9o8W17nSnSurGHhm31o94vMT82S4pD4Qr
yQyNOraFKoD15HJzdtwNdXXNroF6I25J/fIcM3uQJdOIj3jIyO5PNT/0kqtVmS1S
pFwOvXiwchEry8KMIWiFSUtnL63L1ILTMkyHaikoSNpqZykf3hXEIsiEvjTAYmHB
1XlDFpWG4manp82orpyh08jIOxSqWFqnRtvIH9Hvr4J41q3XZHMB8xH421tvIXJb
H6Ll7kIteC6S/5ijtRpWxJ0KmXx9KiL+JlKwmWTS/ZHVRv7L8XO+c8lPLt4Rj+dp
IBLxaXyAjnUwLeaw8qiCsQDJ4LbpoJ/nohIrNyRoXC0Rg/KWW3tkDFWZGAM1XMEl
vrVx2PT1kBMzkBiN3rvvafPCG4tbiJl5MoyM2uYf7EZUB8iYzQU0ogefQXVrASNc
99ckdKyzmvdyxip0nLHq5pv0EzT9Egr+xtmgskRq63InXtTR1UJL5qtgw7RCsUG+
N3dsSBsbYq4iA/7yucTG6muEalt9PYzwitVCgv1lGRfy6NTt+7KJnhAJ5plQKUcp
s5ObvLgYwwbl5cvtVnM8foi7/w3hT2yqqMaza8F0fRzCvHo/Epu+HMHJU9AfUH9I
UZf1hqW5I+dLJHCwJMV/2cvw/A4TojZPBwGMixVoRZNsEQFSV17IS1aEZZrSXX1Z
tY2bTlG3S+LeXsBd8qWNZ0ESsiOyeXwiZ2yUdYyViTdckHgxVaBB1/CchoPF2aGR
WfkX4q1DExufKMVmeRbpL7M5x/k0lZgUtk3KhsupLNXKF5rERjwlNGehYvFmieTd
VFGpx8ZXXiekmhlP8UhUICIylhj/VtVQhuCDx2kqBdMhNdN+4luqzhlhJl0H93/+
8iOmKUOwpifELUtW7tBJ3NefJtN47va5ohsr7aZuNUOrFKEuuhiV2AANTkZC4uwf
m4Lq5RITDdb+pBnMX4xA9usbC06piyb5yUGkLmISlMUxmLKBZTYVn6mt4F3p2iLI
88dF70ihclLNZnSnUgMrbcUysQKum1bEWruuBRRnMQxMRjoKmPZIIAfFKmnyz27N
hjPZDNNaKXLzrarAC+LaHXQZf12HVdL4iAsowHO+tpbEgxQGxmGAyd2ZmyEMXSWn
qspuaTZuSCMKHePXPz/u4Y5LDY60Ni88BPoIj3NaLkl1A8M4MCn6u08VSx/Vhrmk
/MZ+gcIJYu1L1ZGSDQmJa7rkZU0BjA/zssN/LRBsYbX2yqckuK2oWFpfeyt3Hn0I
NJ+XQYxSbwXA0HEloVnvIPY/BLJKiB/CheOC9hU4MO4BngJE059yvYnbJmyXcKbj
kjNdVH8/xfnjgI70Y21TVYQT8UlkYj+gmjPRkwnYsJ3Qi8JEkcEMpTuhiiJb5nz6
XaoK9bUbQPnx+c9xXVLT7L4l+U07r/vbLY9F11fTn/eRRsHxVCUefriqlKLmnQQd
tHeRXCs7kRcCqI9FPhp6oGDUEgk14dzSe89a+P+oQzyWRIG+92qhcDL0YWD9mJ/E
1eRRQ5hwY9eW/R1bryHQk7qqJ5a9MuE+JL8mNmc+Yam3iDYfLHgplA6vfIoEjg8b
6Cpf7oeHOzH7+p3+GGpyVVFSNw/G9CJ1OIkV02EOzb5kdoxidlpSJCB3xhJwTDuo
aHB2jHHFtY+jqZ/Q67qkeKXDbNdzjTh0bQlewfG1g4H6ywLQuOE1+xMTtdC3hAjB
eM1xdfK6doBqtwDJi/42/yeZRTA0ooKV9H5flxfyKHN6cNnfC103Lq2+ldKd7tP5
aVzspyFVUzOpdWmQZl/RCFwy5TZI2UjqotuFBK1xgFL1VFW7XC1SHhiZ1YVl/kPI
YYO3N3zRWzhplP25fsXBxtZ8IdnZfy0RgqYJQAaUy62ab3H5jZcM2qORXLU4wmzS
oWYjgEq07wSpvZ0oC1tQ163Lb2E1D3oLXBNBKB+khfBz4sT1RtGsJYCDL27Hr2s8
x1xq14u2vX+NJbHfcdgp2m/rNzXbWbNlIWGCSGxMAPcgoh3UJT5TZDGF8mBkSumT
f4NHQ/E3MDiMQVqb6rt4HP2hnvkCKYJCmzcu4jMVbVS6Z7VuxS1KWwtHIFNkdClO
w3HkBzAoOcc8S5xNGYJH9TeFM0LxGJHXcdFHion7FrvLbOlqlZJTeuM8wxUBrEvm
c3im3WYNpqtlY+JwRwG21zxNoiF8J6JC3MMudj/AsaA+AqD28i0N6TXMgUhSbcSW
kx/51Pm8WYRMBwMhIc5+GVC/riJV9MUGbgCxTyOeDvkdQuk6An53iNZeFUONA9EE
jA3y5+P/yguo0pcYGqy19MXPyGhBua2ail04nZtoOMiBkMswGSZkALD6GbBKVZ6h
qph2sl2dHLSTAKKkH762jvM7i+ziwjhW3UzJ4o05kJdmZM5p+jZCufuplWRkgI2G
5bc3rGNwT4+Y21/odLSdKv+sbS6duBt3D21uqU5o0uuzFoIYbNDzyx+h/tYMS+B0
EzGfBBYNfvAVz+F4rhmqUYwsNOVAMUFDWnWvZh4KxIdk73EmlMLM6qSzfwjQhtjL
sSO/i/yK8qWNczs2H72Amr3ZLGz01h6bPh11AX/Aefs1DdajMp0yh2yB+jS6D5AU
0kqKfmVYd/xIEuRFjkO3nnjtewKVk6BOX3tTXPu1E2jkIIFWhgWAh5XA+TwcB1nR
eVtnoMpyfMUnZ7VJJIcowITPIRHayy/kux7tnYsZf1AiXu1Y8NZTrms74oNh0uOs
Sa9jGFadDM4WxMNqipEuLit4UzPUbifMlJjGt+MTFjUw4AUyPC/SjeeeZe5a+a2f
kouzQ4zQh1IdwSe5nzUHe/R3BDV96nlGD65YTAmEAq7TS/pyZoosI3to+tashKlk
a1JjrRHo8bDUD/1+LG6xgh9swyqpEQjDGv/+EH0Gwv/aL8nFoNGRrt/MDQUR/0Rd
PPpKwxq+GCCV1gmy+r4dCMxYdOBKorOLpSp3z+7WXC420tNlQXZUSIAfdGVwQUFG
J8Ot9jrEuE5LhfA0GR7Yb5gqGl+WvVFD9jAV3VFe5jZL3las+X804bRbFxvyhHT6
Dniz5Vr1wpE5J/N5r4n+s82YXZpg01Kqysmmt3zfdwFzxRtobCWyP73csgjM6Sle
kKfkAMEer87rYRu1rAKWJVfjGpKzTs0epkLFKH1iUoKFDmKk93BCGD8M2d0vr3Kj
OIe0iaKhK8+2VzKZI71n7ernUh869//aeF4ptPXNsbHOU3ba2ZYTyoXsVW8a4IhB
ew4voiMVWNGXWhg3NbgD7m9OAtBUqJ2Dqpw8a7ejJX0fXte624AsMRmUxgVIPkKW
3E117My9lm1myFtlOvlBgZXCLzg9kZR7kwa/Lzy7JBib583jZ0WSwoj2jLIbwsM0
uPsofSRE37Ft7iepBS1b5Ajbtu9jcwiKoh4oI4aoUKqP16OlCv2LNz+NhO5MaBCE
HTLJ6zrhAOsBNka1YOoKpvk1TW0tVwomcgYEy4J8eVZYIKJzLpCi/HnCukjwQ6JP
N8IMd1bUScajiKAX6he4sZ8fdbM55N9haoWmlfrpPgV3oqlhWpjPYQujfCK6+38J
pJS+/KKwB56eiIQHI3zqFBP4X1fffi1HNAbFTjTDwZH0PhqcOFwctE2uR8yCSIeC
F53X831TL+BXC2+l0WxbGTt5TFfFXYEnLT9ADYyxoW+ijyR8/DDxcX0smBhYo6fW
ineen7yVup1qL5chPDiFJ1tITutmKxBiGu5a0VOCzlucyp/iPqThdC18582SbB6I
aCMwOFJGy3CqN1vBdSnE6S3hrzMZWxHlkiXgN50ItjBuzngQ2jwEoSNz5ybP6h5V
k4T5tgKUzG/g4Tv/A4EcTkBiy9F1dJG4L3kyBktTYck+kAJNZIk65D/Qre1ZbAXc
nGVKock0jx3oAtdvK9BwLMfVGdB+bZL3AQdYmeadR0MfILf8gPh6kZloQ1IYeG3m
arfZw+OgfkpD6cjpmjdVqogFnWTdBEPNtNCbMiK+fu2uTp45+oJXkrRKlLoHEGGa
sRgPU9y3NVHRDpmLirfjyKucOR+uYscBOT4wBxDoYamnzEIAdCQ8rycrzuQHaGo0
mEnWcFCm2HBO4hs0I+N39h2blNwg9cx5y+FlI1CSOGLlu3giTdRPUZyq0Ght323l
y9HX2fS7KsrrrA9xfKlbuW45+MfIlBLPnXtZjB3niayBcsn6F4nk4LWpy42xVblf
GTlqD7IpF3shtsYdssJArgJaMxEedHkA0GsjnhaeAKTxNqLhagjWhgEnTZrN/ZMG
W0DjSCTPQXQtkd5NF7/CAUtH1+4sAwQPJNZNQVBeN4omPrLGrbHwhIWPiLIzHFcK
J7rk6HJaLZ5qGdvmT77Ywl/Tkc8Qf7s0r5pmL49kmWMD3ZhSYLOl4MLnDlkMZznA
/FPpse9g7TbHCRQ/EJevzzSbKF/iuLreXAvo+ZlZ0AwoFdNRGuaUjxYzlYSbT4jw
7Dy74UHTcJWvhnn/aYw2kxUmvuvpSXSMk9st+zlSd4WlqKAgQORBq6Eh12s4d20I
aZkPVnDSmL89uCh7W8iY9ijw0HISJ0PXM4guXeOITzH+aPulKKNX7fq6R5TUZil6
RoPKD/uOegWPdDSBa3o9e+iK7KHvb+pMMwtPwLhA5RT3NlY3diRRsXbPxIYmlyZQ
eAjmo38nAQLZXFk6XSAngpEEpfpYM6FraoOsUlpCuyfsrA3AbTV1nQbkGASP0qZZ
1SoIOrxnEvWkqwmYRhMbQihDhkpRkvy+id8bAuu9qKF/Ty5hlMWs5cJXPyF/WAej
taN7GgNR6AiN7FMJiB50p/mUf+FHTTOioHSQhuwkeX961uWumnH3iG72PEFUR0Fl
uBGFksl+Sajkdz0SrgxGhmqtUePI4qonyybaSIAHIlPQdJrYDCntsitK+C4CqmDS
CYlFry3fqcMXt56u+rI5XvnLzJvAzjfpEiqxcApN1QL0MupJULMINTGFZTSZ3WNM
DaiGRnAQ5LShpbnkDea012F2Plo3Ae15Q58JbyS51AhjAJukBxHRi15RjU08Pj8f
3i2H1vhVnNi4HPGUqBolJ7V1RLMq0yMxbN8ooUCG4k/0V9tMj1DopXeoORRMgnhY
s2KWOu4mXdZTOuNQAdO3m6zbvj0bkpC2BCNoj17tn+UEeVsdn9XjMbziP3UiYE5d
vnxgtSha/2DDJHQ8W0bzq+le9l3QajqT826slODL8XOYgLSv/feRKzJBiTJWhmth
1Dq28/PdyoPmAwn7f+iW3bs5EMvImB2CvhU3SOJt80jbXeBK8KQgCUp1/FpEH/FF
J3dbil4T4+T7jE+ZfxpejPsQT/kbpt9PSkUoV2HSb1thxCxTZS+wtbzFYq8rruBg
ISsGN2VDzJSIJQ80OhqDAaGsbMUCuQ9I9+wCT8RBMsE3+PpYpK+weWJywRHDzrNC
lX7FYcm/crxvHEZ54i9jxl0Y9bC7dqr9DLwWebzQK6rABPhk0ze2kz9P0ISL8XbH
oE6k/TzYUMBOCDL2crGeEJEPcz1hX90wmC1CrZuSoiW8NHAo2k3KdolNOOWnGM6h
HFf9BBwlqbkm4bRaju/5LaWRw5IZTYYz1S+FEzgxo1yNj3vVVR0WpR6Ey3Mv0KmJ
tTS05BmdW4P5fe6vikOwGLt1a9IkxjtR/IUVdWIVEql2adGWRDOO4VxR8Lv+c7RN
/2VH25De3WzHRdENz0XWMINUxnk4WGNLc5kN4j7CaBsgYf/eotKQ27JRCFtrdEdv
ERL7q0eWEzTcrf1M6vEXg8eExOMo+jgfmwLT5iXpYxx10kpjheCLAujfSpigJfSr
FvISNyzlS/7qyEdxJpBJXv3TMtGOnRrKOyqccyeyocwYcWHBW4lDgIOwaIFgk5WM
EviSqaH8pHfCn3T5J87OEbIOqmFo92C+NsqwYcduoAWuvunNEeffkIUKSccQFMZh
kX23zEi0c91mnnye862qci1aVBs4DZbPc3TWBmTP3xTqaHFqsbJz0qmqPeUi5Ifs
+V4azIBXLD2kM1a4pOOAuxQ6eBkrIdtuuB+1qcSIZ90ERiqRmqqjb3H0YrzCaDFI
19cA2JTBMHwszH7LjHhJohMPQWb1Rq6odg92HfH4yuBmhj7m8r3kpsdXNJzoYByH
L6nhLIoVcJKD1M+aDkWGxJAtrU41Sk19F4Cut2NBeJB9q+uZnIXly/fEG10aFaAS
bOOaKeHCeirVeFv9EamQmw8gP2LqmmYhmmXAX8wVzhWYkBFxeeAZNHs6u/G6sXrg
O+Xp1urzkvkkJSSF7In1MJGH7wRjmbl5IByXLfdv3CJPzlsyDB3RAGJO5etdMOF+
h8+Vubz+Qtv/5rSDTftp/CRMhj7Avo/CB8ctjsfn0h6aLy+yYRbh68t4gsA5LmEu
fmO7/TIWcpReJggQ6hYsJUgRTapwCsv0EjsrwJRjL4EZf+6epTGa3cWZyCZI4rbX
+qQ+4GdyYF3Whb8gm2PmRbb8KVN+GARnETL/px+I+X8eL2EKkS5ZAT/g9mya4AQn
ZXnert8JgTJMpY3eAGB8znplLZz0EBd2mrRdFMR63ZTZo0r04rPDyXg6v9giA9Kl
t8N0MlY0DarR5X9EdQWxm+VP3BmjyTABb3l/hwnMKv0tUjYP9k9TeWvgZNtVj94V
N5O9Ndol42ZHkzTxtWRwj0QXZFSw8X+C5HCrpkH3aGQe1mxvBZOGVlVNl5a2KKzi
kPYVyV6qV3WsOmSY9lLfhibQkD0NlA4rW2CVy/X/7K9CZaqr/P370kpnG+B5ZRhj
nh00uWUyObr5kpsCwZYeUJewmsgZ0iLCfuZnAIiEqatKLShHE+JL5SWMAPSMkXuT
fD2dIysD5WnKqBglB7J7zp9PcAyKZRHgAijHV2lIzozubLh+fc5xo0MuGMgMpeKg
EeM1+Tmg0j0aT5fON5bjvIVA7c0x1BnSPrIhbcoo2wOhO0ESqpDVJ9jUvHPBvDDo
xj/1sHWJKIBpdS6KZBqtTwc0CVwZSjX+7WRSkLn9SRO8scFElXclHMGosvhK65gL
N47fITfz7m9xP1f6VSWlCaMXsSCnZquovkF8BWtcjIOwYAPpbSd9t+Y2eDw0G1tW
iBxr7vv0rxma2XFk5ZvHzIX73F2juqH5d++tfHfrcN0cIGT5fL7OB40IIMfIdc34
mwv0tnWwQS0WbM3nkQZXHIBeDmwjxY+HQ0Xa+/2qerrF+5aHBJyvG/Fbiqh7v+Tm
q0JzYsEE5u/FMPiKuIyOQLePHEAdUSyUAx7nu7SgTUX0ru09z4812HlpJs/3Y2lM
O1oKbcQi0nPEvKwi8Yt6apGAO/JuptrnCYXs0cS0dJuH/YJfB+vsmxkI7oiVlPaX
vEv/booFZbI+DaVMHnWOmUfu7YrYPGkoLGldStw3CLIvBiWoHRlW812vggkpsDsy
jAf2oZg2T6r5mfYDRznKTV5Rm9T7sQq02KrbSgWMKioNEjdDwuXDf6p3hX3en/8R
DA37Rw4jAc9eVTYg7wFKYyg/7sfOaaUFNsCM5xFQuzJZQbuJ78+szltKGsWx3k+c
D7Rs+E3pJEj6UlL36nCYw6MWDHwpMoQ9FA0VHqc2tT1GtHQXjSzKEKrSe+6R55Rf
qU7+fY8tXOeZdRPWoC418V0HOtHPlspZyAyRe23XS2R0amW9iQ1eCGOBPZXhBZEo
QUZYOmSat7FsPkZJRQliW3XzDL6hztRXpm9Zf/mjt/8CbODFtmVxOMKOcHMcFLKo
mfAVGsXzR3Raa3w/RyBwEZWKnTb8aeof6eDc8ujzbUJyqPtXgMFXO6fbxWjTKHBI
CQRBJk5G/z5yHJZ2yTph87ewjyzUOxvnVmWvVNOu6pRKGPlbV12oUGkmGaMYqF2B
t005TSCTGrLEj6POzD+/tloTAkFONJJ8PeG7NpxekWBsDStkRGgCSshZHpCVA+iY
4yv1L7jm2Omn8Ucu4xOZpzfvPJap3Gw4O938bGGaZmNllHWqkYNymw5s8941uRsV
KZfeXhZbQy/IwjCWirNi4oYlv8y1eHP2CnxhfUutahECRSo9y2INiLIJSs+SeFfQ
Lf/2AMYDHafo/0Kq65KkrnFC0VtD9rfIa7VafDeadELuNMmAVWGSR79hdyn4MjZ/
tAcKjqPmJBL3vHDob2L06S8V2jhtNv/iC+n63+j47WRIis5at8pNwNCRFM6+Ner6
wDeaHfeuS6phm3HuuiQ6nBmehtDmGIOk6bie/+8rZQZgic4WEpFAIPh/6ScHotEn
iSktLUX2zq1tB3L9Av1lW/VFPt3jNPBo9bme1UQVNeF7oWucGaklcdOUwywskvx1
sQPC2o7XSFPShnbmZ/DzrOp9XRj6/Zg6bomavqnS/6UeQrcTxsIgf6EiHhiWaDlR
0LpfkoJQHvhXNNXCvBYvAF4SQqVwow3x0hCZuh9w8tpTEddW3rE1vhzaUKUFQD/4
0EDPqlOzGDi8SsAUr6FUsQClLN4ckVit8ghIzZGw8EPAeuIkz/STAi26ZAYE/6XO
VvNN+dsCjsndKpRErbNYXmckWvM3hO2x41gATW6splq0fUgWuZF61LWdtqfjFmBy
3QHw/bWmAWXraAHVONHLSOgdpdSKGmeMrsb13BlDAT9hl3LYX0Iff4CIAuvFvFPH
kleguAU3nQJ1paGQ6TNpwhHHkbWW1sZZ6ilCP92/j4YUHTaRY52CnbA9LLXmne8G
535SgZVOIjMqA55EkzyOJdZIXzeSQPuEfmd0A7GYzJZ/VE6pu1hXHQkuN6XORzml
LSfOsBiHZvBkBFAk9NgyVvDI7aqbvI4UJ0HRvblqBOTGbjJCeUCcuJNuk+9+Z9lq
dTyaHXHznaOJsishLZk2BhYOrbt7qQS/wbwMSwKErtbY086zI+r/xA12+6QItRqN
idKDaoDjRp3est33sJWnjC5VwvjmsXwlO7jxNH8v57DPKG8inbO3mkH13YRBhoU4
b5eg52AlKAspIvBcEUhIlrar+yAD5Sz6tXSZ4ORMwT5ZLHOQ4SimK6UoWqAAmg8U
Xe907EK04w5i4r3p6AGURL3ALRCDSgJRRKVRBXgM2JTfI/5/5TE52hq0oazcZRyc
Pdd++0XjldIMEShdFlCAHSlPTy7nW4SduVc1qafKg6zFeknMrYVnlb/OFpSgvGLc
ed3TsLy9mc1lsCPEZs9VyW3N/szyWuZto98XINvhhsAm4fD9ovbgQq32LNs5X1C7
hTV/z7cAQob4rJb/Vg6bzr3gw4zWo8Q2+xlWHUSbTkzwGVowW7IgYz0fp4jIhCjy
d+gJfNzjlLT5s+WtET+y5gtipq5KVAkrSez5W2StQKQ8ZVrGMmOZCCQSceu36FYU
5/HhzXC1ySyfvdp4WA9O+H7CfbPb5FSxwT7wJxmaIc+Hj5pHpV6ZK2kP9/aPs/eG
RaIhASZaYWwSjN2zZrfAqqdZ7x3No5V9rYroQdJjJaZr+HBagODO5T37DpQR7KoG
Y6qeSrkQlB9fDvI0Uaod7RCAECF6mBXlKPlUBRP1aQgSp2j0j+gQZwQqsD2fAJYJ
`pragma protect end_protected
