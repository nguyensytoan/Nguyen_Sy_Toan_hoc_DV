// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
o3V+hOHJsngohrw2TKOp1XOGwDUhfpOB+ns3PDR+rivmFT3QFGd0W1bMvE+KWQiK1bQcsQaAMHXy
26EqdYylYKPwJA6MUlhZxNoHrU6j9V5Z+0XZEnoPs490CmGOE4FZOYqfZU9dwNCbmPL7PuyaWStC
V2ZdMR8kn9oddCDeA+f7+qDR1iZ9Wj7EmLV0ac+dpye+h+hn5LLHG7VsDOrMT67B8XyaWMh3fL8J
s+dog6T2azrZZ3jZ9HQogTKI4l+N/MkIEMA1rojzIQBlV26JvI6KMHxwfkPfeNAZwdVA/ZAN7HwE
vxRCpm5nDG9P7FO4kzrUuP5lhtM08fmVgSD4vQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 48864)
WlP5eX/Lc01Vd/hS0v7Cosz5YK1QmCfseRkjWSVmutnSvE8RDI1a74F3r1l0wc5D2Jibm3v/zl7F
DW/c9yhaNHnZhdyCDqN/N4gssPylRgPl/nb0nEzjcYWJf5FmGbNaehA9g3fbWxKDCJzVVjQP7B5C
/quxaiqFF2FmXfEwwQGxxnheS1/ozTW7PVTAlGgbgBw28NPO3t6yOHW79O7uRkjrTVM5WLAc+Ad+
Arm+u5NFjJ8fRxV0MOwyK6uY/213z0nmM6y9K87ofndH/bmLTMLQZjft7T8dyJBDMJJhz/YSyrsm
cFddQ3CChccWrYE9/ompz5TISR9bIjptHZUekRDGmygAlkZcamRkpK+YnCgu9cj8PO7bbQ3cOZiK
HMSxf/OstVVjgygPeFWVc7dkcD08w5BNcRmQgQobt2R1eMnIdGPXmvoo85ScTuPk0MFF/eGZf11W
4AMDEwuG6vQV8TQEEnyUAh8OBASYSoE9n+TVwCIEs3/oPqJE9Kbn2i+uGxaAB8myfy8DHNosIsyf
dX1bGXNhrmimt2LO2qJx9EgXaiRl9vgyigWZopwRF9Yt0y/nWDnORnprpIANbQTDB3K+jElKNTtZ
ney6FeQasw1xzEGqGuRWbRwzkPgWJEtIZqjFo5bkOAZTDOtE4F7kYR3n6ZMmaBLFeOoVzeRIiLaB
Yq2iboHpzEQwLjVQ/guJcAkzfVapyThPiH6bYwV4PehauIdKXbOSZkimB7f/F3ryCCvO8LCo0UG5
E8pzFQzrFrD0hZYEC6inR1kZcq14FY5xqsykndOL+Z4oIDgW3fZqQ9KNwHEkw2wiCbptykLAROoy
XTYuUJyGIqnS274Cpwfz8yECzACn0amD6+nen7zpWZV8g4xx5SQe+H1qzroHfTwHBQnWMY7IYSSa
qIVcur0dpOW8ZRSYrUmn30TTwNbkCHeiwZ3Fi8TlQzKKUMpeEfJzyrN0t02eJhaIYSif0dpn+DAe
wUuH8PRA//68A7UdjAZPy+u1QRh8v1lUKW5Ib3smwbepyPlBj3Wjxu1tTY9yUi6b0/h0ytPmkGT4
gHrJsqH2k7SZXhzjtlZR0QABUaG//T9IdlJG7UlLnJAgkWXYOGNcrYloPXY/r85WHqljAfnUAKor
TtdZYD5c+9qeR78mBkrLminvjpJxOk4h8QSkjGxx++4lbnLQsXy7UXbpThvKCfWzgb11GZQpyZFj
RadUS2O1l47DjDxq+HrVFMyfbAhwbRBefZHD51/1gMpdFZYgxQS7FlehnrXII1XzCLNrOnBHd61t
TPJ5yK/c0yX/38eslFc2pOpGpIvYcAsDrNbDTBBXNudotIEX6M0jfYU+WgP1ClJEF3zqm47ROmzS
sK1B6LcY4Z1j5v6VttJcMFRCfWzOkRpjr0sKSmcThN2bQORzSjxLqfpuoril73zr0/A16kPpNuNj
6nVkWEkExLGSz2ZLz5zTWeO1PbfugGxVLkvuggyV40ZTxNdapb/7P+jwT3Tw78TNNnJv27mkdFkH
cLaaO/LQ9mIZzXfEChb0N259Xl5zFcwksVoikWhcOoCNq++Dj2X+5UxHWBaJfhdK8k31/7oH0pUW
G9EjfT6SR21qtVfr/ZDIkCB7XWnAUMmb1LaAyVLXpaITzOnHQ2km3tZKIp5Inf2ityE+znksUxPz
bUoiOn4PWgjk5KA4XdJVjGgxnedHqb9JhjlFP+U8D37r7nLbS5tkJjDX5a7Ns7dcgMaBMsBGzw2x
QVSDa7aEFcNa6xDG6mCWzPkDlPEFGS8FZlEpGm/SuP37JYFXAYD5lPmXHBsw5N4+KILQdlLEE0F9
pL3gJ0rU0FJ80b/10s90U/w5SaGqgWTjOXrmMq6wpGvUwyC4AzPgqKBc/lIM4E3OPJQsoDnS+k14
Hqp1ysZGqWD77KsyeYo8RnPbC5lnFWhaPhST49IbK1/45IiqgVmMRrrCvBIgd4DDCSxDY1U7sr1j
WMvUeWy5h4GjIUjz+4IiwjTb9IGWdQC2mbtp+0rH7CUtxTkP4fwbxRcO/aBl7f7DRiOV44qUXQVb
6hnapOkBWVNjG1LRplDJYQhtypsyfkoH3WvBZABHfZwP241zM5s9q6ErZDbfkQWDCndUmNwW/H9g
3+o1lp9h2SnwfNmIeQPavgnT43u9y7AXJDPalv6bHN+789fmRb8kCkCMzNKdb9BmYNKYZfKuahwH
cIOC4kymnF9Y9hmMwME8bjzFlhHoCcGnbWaqAGD4+uJy6tgXUZUr2ifb6MJWN3HFhln5b2vwwiYn
kQy0ABGWH3DDnjh+awqvuq5VsTcrmDDwBkOkldSjMXxXGzAXfOoxAzeThnkXJM0D9NTytaUczc4k
qsSrVNBXJ262rKVzTvd9IHOuh6r6jhZa54svVcn0RI326Z6H2Ek+2d7jswl6ugBLfj3Tsx2C52CE
yWOHwgEtH678KDycKp5fOy9MKPhoAJhG35aMyhEYJjaFJaxR79fFODG93gzXHRZDjmuUbcSiExQw
B/dqqxv6KbNURQUHRVPHCCf6QiAeWBijicvpJhSbKoSeqVrpu6r/oMsncjAw6VQSIbrX686ifdZw
h75hB9tDfxL8dW5VEnhTe3kNHzZUk1dbHpkSrllY41VWrFZZEHzXqMJ12mTMTs6XNwpIv44WGWWE
VnScN6MsGkQjcXTFG1IZ3rnBXL/5PaOEsYOiVnyo40Fs+I1Jy3WxkoarTDYrpADZw/x6eW74v/ls
eRz6lG/Rj3umv9C3hae3p+XqBtgnuw21nu0TPWSTbdswDcGPDURwsOkAO+cuGLgxipioPyRvRdix
yNh2qRUFAZP0WnXDZnU+/dq6BU/gBdoRLfXoaNBChp0O9g6WY5lUuDQY/iZrg2j+ElnDQAKbxK0i
FbOhBMJxU+Z1+6lNCEm+XoICQD+79jNeV89nCc469Gz/N/vRWXgD0HaBrGJ07c/n/Pph9QUy7xeO
Zf8bnAAr01OvcQPQaDlP6d+Y8D+bKyqbn6Kag4OuOwaIk8/YzLOwDWTd4UomoXHF3/2RARviE62p
1wRL9P1gs3K7OC6f/mtlWrzaYIj7ZjueecfofwGxZE1/h578IJs3w2QLr4PNrdEKvd651swlI37f
3IRc6G2mLyYBF9Hg9giOB6TpJW/hA7qU1taxAQE79iWcE+HFYu4Tbh94DfEI9YV9iT8qYR5PGren
75UFk66QhtGVhJDY/K/wQ8lxRqX0wXtsm7CKzIGmEIZBFdKe5vJJzQnnW2j+tBK0Vy0qCSmdisE1
54q2+KSRkYuZ2nU2IRY6gdCRo+Kl6hPLUXZmMOWdtopkSNki5owp9DTLtJaFpEns/NW1GxzWYPKQ
xAV0OauSGp+jZQJX08zi3WgeJkwyo5TLrtl2yaha025FLSzfsdmd06abmldxLIdKxk+EquBZJOuj
K4WYWyHZTfGAlMxGCVqCYepuzPzQQ3acqQWfNBibbvMO9SJAxxmwMENke/nA6yUB+AvRkkgR/lQ3
AVeHS7IWaTDqwaZrbx4c7kdIiC6zpaWC9WgtZC0cPZMq3sUq2XpZXHwvn6eWkXL9jNNUaG7vXY54
5JHljEK91rsSQTnW8zRzNp8HL9hVxQ+yKEW2YCst+Qee163R+IvyoDd6APPNCIT0bit6rQWqXiAY
SdCEQcChfZTVgQNw1DAmpm5v4WhyHXWDCbefiHepL/QYS9EyjgvhfqDOogEvIQCV/lkD+ezafDkY
RZPCAywpsLfijUZfr2dQlYBKdOFWbMlskg7pMXIb1mUQ7hOZlq5XScSS6F0NGK6e+ddk0In2Knz1
HCelADXSLmUA+jNvc0K6IRFkWqGxaK+S8YjCf8f6v+w4VzGxFWKeqXGVaquofQ8JeAziqS28hntk
TUoURSpKeNndu3qUy6+tO9RfzFDMdEfIP3NbRz+t/Epmv0dyPE11KgQRrVNJKUF/2foRmZR0ccGt
YY+1Ct1bUjVMnUPLwfjdiffCTgQ5RmnATcqwCo7hHGEH9OXEOL+M4aiow1h4sTX23sGHE4OvvDJn
ViZHWWJm4+d49sKWjdNFvdc9Kja/He5DMieJIdwLrqy9s0CHSA52RhGvRf0ZN8bd/ZYqrVln/o2Q
dUIgyaBZG1I1ReED3fWru9GCNdlmn1RgBN0HG+VrtJuKjoWwLQIspe6vBMNLChKQv886mFWcqLo3
S+Z3HoE3I1ZYFJ3Qq5DntF5kg9jB/EJSBiqun/gd0Tg7RjCfXR6EFsfC1Rjv36qUjIdzOlsXpvoz
6XSijASFOg+seC0CmFkNpigN4KG9sRFIh8bFU/BPzgKcBLkl6WM94VV7ESN20CbNH5RP11/GdaPt
PhDWl61XKhR39Zv+6Yc5r2mt9p7HQhJB9vWAVZTVd265cWamF+P7KkeXTfFHIZFRWxUG4QAvk9aU
8plMF+FfuKb4n5eovGs1ggXctXbMmGO/EoxY39ktKAwsAQe13Ld2LS0YbCB9LuNMu+fPU1OlH0+l
CepJdJk2PR5H8mozwZ81x9/7gJ6H6pE8JAhYRXL+Y6jT2qZ/qCjaQN7HWbFVrbLNJyzX3sac230v
LOLXZBd5HLbvlkp1ktHJIGKSeOC/E7y/fxSgo5iY0/KIcx81V751XfEWfVZagZiyOKgIZiOajjkc
L46FIZYoq7PCcmGa8CXeb/+l//VZpOOjRsFEZYSaEgxCzGm33CZLk5CXUqhoC18M0I0FFVSi0kUW
bBTYIBvdN0FMDlpu2YlKAzPWFerP09hZGnLa6xWjFBA4YJXvBPxjMIV2w8G4gRtKITq+52KA0axq
9PIvmbIazfDz07ZHrhLfhetL43CgDplwXMswZCL4pwLokOdeLHc6aUAunztmtx8dym0iEbdIbeN0
650We7iwB33Lfwl9tS6VN4Z2Uk1npsQ3iNy0p780J/l9wUEQE0rZg/8zzzD5k58kjAX50aNb4VNi
UaM+hbZbgHAcQeEhPaUZK288wTD9jNiTVtLpvpSSBsSMqoXLZw42y2RaJsCjZ2IWX8AgoVO+ZHox
Oknv/AXJIGI0pBdcqLZsT33S1src4otsTK1EImvk6MuCsS6KTRSeWnNt7Z1Yd6WH6TbEX2tdN16O
tpE71E2AIS2eUsY1rXVnqoqojmGUzREThQQh9S0tfncvCF14SNhI5FQ82fLVsHFPAN/vAyHRaqi0
9lm1yFQ3YZGDPG14pi/qVCXE517hXrz9zf2oTmp3/yFYfEu2XJxc0jrM6BOZ9piejeu1kSAEbJy7
qqPUpaoIciyg/0F5l5UbQbq+6G4fzZdyxxBeSPk+EGFX2UUYKqSdJIdQPw7ac0naou/FQH0Z3c8q
8gvB5V8LY+hkOU71atWv8A0SJv9fJMRyiCwnIqd9PCUlHt++45Ezrjt2mIdfQt8azJ+mqJeKzbQq
CRdkHMsmiPjAUtNaI1axWlNCqLgQz7RiQQAstEi+RzPKq42jcRjgLQunzHgqLQHEwN2/hwByvfhJ
PuOqXZEsiNxhA0vWGKygvHB7580Y4U390BmUus/xs6rXRbIvMkC/IRNyyzng5gD+RCmIT7gn7ZOm
dZuM3xAfBI4niJvqJuJO2mU0JDYlaKo6tp8Pxl612B4xSJr14QnGi2Y/NdYycCmwrsXgCdgVqxhu
4mT4pRfjRm8Plxl22tLhF75CmaNlBRfFbqLNqHbFbG2CQgPHthV76ua011p6NnFcaOpnPngy7P48
y5zSzYpJB9CA1ouWHb1vW+CPZaLs1yOrqESHXitRmfgT4LIbm+LsBV1lALRyeEfOTte9/aqXoaba
g3JfyvTcCBhyJUDw5lS1M0DRP7hGpMFvWrUP+qhlQ/bDl1JKqIv4Em6sQqaog2zdaPHqDN0fIhb0
rBXouCcG6FKX/u85jdORkVAjIZWsBNQkB7ZENbdW7dUk2qgZ7GgGejf+rSH1u/hWR91jLoJckPOW
qdcvNGEbKc9Y/PTABpqWfX5BNa23I4/jtwgW/LIBfjxk9L9Dx2bXnK/OdEBGQpvtvXOOluYOBH0Z
hqardXD/AMPjiiImfJIhycMD50zGwEyQRmAtT5zIAKMVJ4WIG/OA/06Onhnq8qtYVgoHpgXK+ph6
UZbCyywys5ClaC7MYgP77g5zzG9IlYSSCMjDmAkjVRkeZ1moA4IlF3vQc47ZPpKuzM0Jumt/7b2S
Nhj5wV+eXOVammvDyirQvbrlkcrHTfAT+JVv1vGUC/7SMdYP5QC9r3R6O3Zl7ovgPjuqA6J5z+Jq
H/hiIZjn7dpvcqH3dyGIGLQIhr2qbXEs0O3maqKO3TpEXG2n4qaD/hYHShHy0NkMDxSO+nex6JTW
vqaLqYk8sTkDJ+pLdCIfBYguyYKFyO5dOmkNonPCtD1FJh7X9cnfWx5QhuAR9DrV5atL6x5qWmFF
SfjPn/C2s/Z5lW7cRKykSxLECzBhX8wInRf950UzeXgDkKz7JY4KLBy3q8ukH16HAKySxtq9lRHa
Gz92IXZaGLUiZ2WcYe8qYe/axtD9VWMmaYcqfbOgwkz7nJAtI99WtUPgIr5mzkPzOltD1lzI0jFg
teDmMoFXPAs587gLM6sP6Gz/C+d00IfvsRPQYga1NHkSITsoHKn6zNg3l3gGKhUocXdO3G9HE74R
0ryuuVzDxGy4HpzJmnsjIy9F8ufr6JPYMlBhYdjeFzcUr5PEAyunQyXau6avxDajNoPWJuKhDT+4
clNpS/CR/cc0WcmwXpNCsR9fBPKMeb1v00Uy77Q+zunighFy5a+Z6fWeVeMlNAK/TnMW6xE39CqV
PcVwqviOErOI/jvf/bHipOD+K9smNfizyrMVyRPUN7e+u6mWY5up8J4JoMljMycMCs9xEVP8CLpn
E3BYMTHSNCKZpfxknYK6/teYrW2sLHdgw3mw6qt1uuAJYbA8G7uwvE7P8BXfOKqgNHdakMJ/KRXZ
x4CvowOIJSwE1ux1DTq77XGOPqL7TFWimDYT/8NtIUYDXKIhY4r2kkO0im2fKN0fxlA+kxtsoaid
vBkeX1dqiNGdbeSHvtXjb/a3ikXRlV8fMBRNvV7fmeEd++nlSlndudrS6cavOX1ev5H7UzjeTyA3
64lc8795I3fMM24U8yvD3ynG0ezQWxXhWQ07M8/VDdkfMxj/YocUDxQiS98SPLU//wXZx9+lYs2l
FD31SN5kSmgnRPWEv0A7z4c6q2uA7Oy1HLFs9mBagqqI2Sk+lT+s1IH4cx/Qfud7z0xkXFWe6OKj
q7DJzIlsPtmjhRAFJ+ejNCfqdzgb62feDLxR4RNknJyqV6Hy83LUysRxr6rpAx28gDJZdN+6HEzu
mCiq/THVdFaxxWuZdWCg9lgqye7muOgIcmnJfJEjAB+g/aQKCYOwAicrWbAzqn5oPDwKz3NinHZN
NqwJVzoLK4gwZX7eUx9UOqPMpKDTvRKKzL+zHr8dbKvz9aMnah129Aqe/9dlcJOvmPYsXRK+tH1P
FRf07oOtmWB13Nj1FkPtYwoTbCItLK7Wf+8qDTwQ1oWB0cojlIEtnB19XMgpmMUUdWe95cZhtgvb
nPEJHBcplmnoteohZ52/nCht2Y2gaC/aAx2jfUIexJA4YBgMqQD5WFJgSRpZwke72KiONdLDDkfs
EsD98ia2wIQjng8c4IwExBZIIYE9d5oUaPksN4i9hW1JHGzz2fTHyHw7Qsy6QZ2v4wmFPoP+yPey
Pe3Uz46dwlRTOANUmsaCATVpBwiQc6SKoKGSEb1kvfRBojdNQ7mN1txFxprQvs9R3KzPEIc0Lpc+
+rg9aU+WLCQpzyPy3UZ28h8fQcgABqeG82w8d50jTY/kCvSHrXjLW3xA+03lFJ/zQNpaDGZmmItJ
7o/Te2izJqUlQjmvtjXBVFIFQ4f+UM7qUTjBKyxmSG99XKTpfLgoo2Z9G1jNmYsloC2gFDMiFG2d
eAiUVavMM4xqEzqtMmQGuo+yaP+HDb0OpthGW8HmoJqtl3y18ovhd+jGQua/BiDxBpHr+w4bL0SJ
cAnlF4xrzfWt0mIFXZ0hOnyqzFg7BLucEcHGkU0Xhro1hN5N8T4/UHZVaZ5zLLIdCTuN20Ded6xh
zVlK1IZVoOVsYk408Z8LwKaLhRoxhfWiDNktTNd3+8jGQGHD9utj//aqbpj0aiBmbVtxbgJKKp2b
QbQhv5/DswQd0RAyc/yyF9F//92SF7NM4Bi6fxkvb08rPSdySuG0RS8wK+CBVUIQCGv95pi5VIWi
kPRspcbXw+BDLfvJasQN/I+ypzAbG9ilgj0+7Q7py/lvaH6wHn7iMRnVtSHxV3TI+0XAfjkk7Smi
xEmnU0MBAJ6QG0yNlm32c6EgbPxeJ+OiDhL13z4x2wXpvf94g2+713IOKw8uojKGo/YNh+W1DFND
Z9M3jDwoCo9unYvCNl9pTF5FRRyVwPRHUSgxvkLGJbcRY+yQXKFR+AC8IwFnM9GW6qp9pM0JBHP/
DuNNj56Ol3vXliMB1kkKYEiV+B5dSlblZBf+j/Q0YPqwniM6zvMgL8rpON++AZy7uM5Ql9DMLwRZ
V74A8zzxUka7zrrk8RRwYmmalQ/O2FdzzyEGfZtj/lWlr47Cbxc3MaDLsyvtfKUAZCZnF8mhgPRe
L8TPhxt+GrJVhgHP5mdp6smZK/VUzw64pZr05+Vbgs/9bt+bI3PXIKhShq7+S3uLN45d0KijnUAp
J+5zXvCSlRSMJOO0rf9nSTA1JueNViZwg/e6Y445iPnAjiXjuqTbm4F8252sYHnhYc1TT6fX0EMS
nWaNTMG7TynKmNimEvdPT2QXSlMe1PUEUEkQd98WE7kGMuT6asSmU0kjhekus2+bT6/+xlUCNNMA
LEvCngVl3tl37v4TsNQTszhqgvPQI1PLgm4E7bJOCRNzWdA8VVk+T119qP/Sol0/DvrHL7t5dtGe
9+I164VLjwGnYbclRXoTCzV/Op+l4Pztw3hs5SwFAjnlsrShYgygXL69IhWL1xe6Ieu0YYb+5O8h
unl1Kq3wMHqAYDgYE4hePxfe/cpMC74FlAmKwB6KZz91v8bvtNv1eLj9Sa8sHrzntou3ateunWUE
BIeusf09PInIigtGcTul6F1/u2Tr9WmehXf+Nara9Y+Hmg+8d/bR3cut+Msf4wAT84GMvnb3ubwd
XEsULxvQcLs3JohF7okND7DvqlljMs/M0BT/B4/h/9UBRC4YEyKPLGyj+K4Oi3stRAQwfDfxRa7I
S98skLr1j3fc3t1uEDqzUcAqJGnOtQQQAOYkKOFUQgvFr8YtvVykoUnqgl5nsRutYdP82kZ9C63s
X85CB3MOXpHCDtbHrUnnIiFOPTFFkddPcILlJmY8+d8Z/fN9XmKXbyRofCw/kyzeYmWuKjXTSByF
NHaoUHa7vVruG3UKFzKoikeY4bEErpgkZJ90+cx+tkXVVSG9pGMaFhSRDnhY3kVg8qX+aF7dEybU
XHOsNHueSgLilPQpWnqUXpm2u7W0kS/cq9OM11mTAPCXuGeaYBk5R9wVfSK/VFAI3W33jirNOv8i
B+4Dk2XM1EflxAyzO2t5SDhC5jQNhauj6Jec3K0G6ArNRnLJDIfBe7Y711demMaAVzI1GtJ1L/OV
Kqg16X7MO4OZJCMpK+gSGEgJHU65PbM52GFjjc2Tss3PoVKZveAyf6L3+NUab/2kfuGrLKGDE7Hq
RpuUD8f5/1LCol/75Fpe5Bs6HiuGKViFybrVjlS2j53zke7cOqas7RmDC4Mk5DzP+5BIDr8YuimD
ZRHnJbNfBrUzgr2fJ94K8f7s5YztDfz+yWQll0WlvfrUSjydQeB0aknyRibCLJyuSckpLN+M7JFF
wJ2Md4UzFcHfdzV8qObHXxoUevmMkYF23u8HY1ApXPp/4Taj1x9PAcvwiNO6y3jrifiRlmeYE2in
ZpasMTOHb9KgPO9yNq2wmDM+DqAX7LKcV+48+LNdFdQVTsz1FP7ZRu8/8KUgBfyyICO3hRWGOZUc
J9pVkM0TmKhKMP4ht3sGpcnkDIlC/W56u9366W9N/FlqqFtCutIQz6ApuXlHG6xW8Nz4reiZxUKe
iUvwYK6eVn52iTeBPzfuRxXvri3+C7Id2P+yyKC/PuTHsKr1SOWFmQkCLmcqO66QM78Yi54xUI1n
zn0TmW/SgUETJJiwoyd4TRt2eMtk3XWvaIOObab0eoTFYCuSb4+U5OcYbnyf/izEzw2H8Pb7xo/T
aOYDyh+++zM7IeEpu9QvZkObZ9UP07iaFgnc1Uk6+0OE/GR/W79OSw9NDkJbw3j4mp2HMZ9fy6qU
AHKaR9JDvPonZtvmowiLup+Guz7VPSKrICel7O7oqCDXlsfUu3h97+MaB+1VSrl7dG745H78fGs4
gr5+zZPR0CpRM1qfvBV3NyhvV7GdygN13PPvzwRN7v0flAL9gSI7OuTcqtALKJtCYOSdxZC7qyxF
ySeQ7AD8hwpZU81F7o8aArvnvco1JFD0JzHz63k5T5FXjMD2hhNfWUNTfNR9B75DGlIfnnR2x0tb
eOxd8HkYD5vCXPUN5n+4l8M17bXzmB9gWpERlTEzUvY8Ain4T4qnvmcb0hNSYHdf5qbrPMo5n625
yGLCrKf4WTRIV4yptAz96XJ8qHvk5bXk13vBAgyg8WNi07svZ1+sr31ERnsr/1ug/6kdQk6uVEvK
INhZqMKmWnS4bR21Oj7avtjtazacuIP+z1MQUaJqfbNQE1D8F8MhyaeHRiL0MFqU4/lV6tX/tOPy
hT9qnwWiu4UC6JqF3uTewiE4LegsT9e7af+2l6QAT0Yv2Bg8ucWLgsSFV4ql7pRab1cFG9c2IeQs
nm5vk3UKZgNc3QSl2CAEwGznuNhJmPGbxn/X4qrLJMvT4Z7wOmlB3WDGGTmazTr0hALVihIz3T1c
GH5OjoIo4L3gfjDtbsZd2YrhlmqHT5K2PatRAKqdz7qHqkswxGN/kS1LqM/laZuxBEOh5dWG5Q1q
zWpiOtvo34sP41PFsJC886qqwEBN/nLTd4TIZiuoBZJ30fOx0Ni+i4ITEhVjI+9eWdDIMOIikuxh
1SEeLutd0qI92HFB1twleKrNBFmtkzsWCTW0c4YdjriTy2MXKGgpqSmpdAr1NxO3UuJmMxc81nqq
KdeGjsKTJ/JUm7F177mfxMxj6u/xbLtFfGfC8EP25EjIXavjsHzFwEu0jubQsgPVbkNi32Ndl8Pr
/640Eu9e5tsQMpx7sEcMbNmJVdst3rDPGzCGkGToczojp0LV/RrTZXhi3fnIQtMhmStYbt5a5tCZ
4BVb2PMCW67LkTpLrnN5N56u5q9CeKTs8L3L+7+ZEZ9JDFNAqKIkDgB3Zw2Y+0pASf6BZyM5Wh9k
jnI0jigBYv1h3zPVakf6scG6pcKOhCGruQIhDqxGmvHWu2l3iDqJk9DneiVyWoOLsX1+z82lO+lY
vmltMZuiL9AJq9eFq+QZouraB6RKLS91RnxvVBN1dBCBY7XLU10Zh+gTqd0QFKDYYYGqMSYKMTDF
x/OHYCkHOKQmxeZ2qdAJt+21H9z4dt4rafGR2zwh/0tWsRI5BZJawNVQJYm1AjSNFNgVvqdZkT2H
QK8igug0wNSD9M6dQlkPQhiia9ooC/rLgXawjTZZJAMvmuEm5VfPXBx2p43DvUJSRrsp+Z5BaJ4M
SKovGIb186ZgYeBE9MoSpaqg/L4r/0cHeinPqqGbItBNoigEGAJhUaAaHfanOaSBliGlRTZtEjpL
BMkEOuuTWvhFDMqCzcnOWhoxOJbaoWa5+3FJFzb8urvVimufU1//4YloAyFbITLDRWqbM8OsYxlh
WqsKMQuNeAes0B3iBp0l2wzZX8HbZrbLdkKBR3tzPoUCHfcX4oZKokKjPTYmE2pfaNzkqFoRFERL
JF8376puMG7GY5GfsXJYujhQqavbY+6Fdbvz3zLA0lSCQku77+9JI/FO5reOfEZmgJs6/06sBrET
e9+b2M43Kb48aIf2f0eYBf+FibA7imVw5+wAckU0ixFkh5zCZE8XrHJYFHPb2BpuaZzwr+WYTO+2
HGxbyiqRcuNAHCdVeaMdrZ1IwpD0iWMI+zFtMIdHfqkvmcDMquaxewMK6/9XPjTludxcyuKwzS9h
KcbvQWEagAvZctf/ovtKTHNk1JJWMvmVmX1bcBpU4wcCw0r9+Swz8yw00u8+nSs0RUYoTIGZNwIK
lLMNXL59gNkwqg65FausftC/qt8+1HziEyXtNWqKZSwHL1/6aukncwLEUMRjWKljeMp8EePR91Vd
0wHtRdege0nM9qttgJTYtsS92wiQhH9TaQhrAdbKF8VfesiWzkFTN4zgUAkiQssPsM9615KjkkgW
Hp4UEQCGSOYoTARdqxTOot3Y1aPDxfyFlfJD9pMUnc9pGcRV/kyTuiU2Scw6R/esRYkmnWgyaApT
gz62ctAev/B2oxbFirGBxry54fUrB6+PwNZzpssQ2s3qo9m6mm9jb/x/p8PWL4yG3kC0+hYt/aCK
UYodQlLB1M6vOtrWxY0ANv6GB7j2PCxjbwaL8Zs/Ncmw2jrylyBWwWrPURBO8GpJoWvYKE3RWQ1C
Js6ngmSBsM2BGW4O6PJ7oxaTqHy+6F/G/zefwI8UEXb82nHj/GidD7ANAGH7EZRaJpEFuBHsN6+D
eK4aQs2k1Q1qBMmA9BkOdbSxNscda32LjxJvTu+KNY16ehDmjRWkVuQp1q21oGIAjCP0dsVduGWM
oHvJg2fS9yMtRUVhisrospvoTQjtj0iLA3ruFCd3se1YvL6gZxCiugLl39e9DrA75o5tYFXbK0PF
CAnb0olfkJhV/qJgCdDSgFYsf7ryK3IfnI/GRcYAQv/ZaRSZe/nCvfrBDDh3bGW7Etd8gfpYXLq6
PSAAFJ8XctX8oGVzJSvy2JulTwszhh7/N31a6FifPSbD6XJpEWZV1h5vAmstLOEEE9a16ZKjXl3h
0eIXRu5qfbKDfCNkjD/yaCd0U/nI29ZVnyRUzuwfhC8uIj3e0OPf1ShEJ/nywvrTKUq1y2NVNrMf
xsGhorQD6Cihv/l2tGOVzRzeZjRQr3doHXr3JWKRhYtmxpsnFPYCKiQ3hus7KiyMSw+zU7KwOcxR
4yKAjThgkUd7kpBhMeHJyvSxJ7BrP4mzv/BzSv3SRWR+O5sCsyIfdW96TBkyKOxNhkGg1+TH0JlI
XmC55PamVGqSrQuQi3KugKbDw0xa6DAosWcDVZpT/iHGfUQKr6Cvm90lpcUK6XCzOrXbyacx37L1
aWaPIXqJSEGnVksx5u7YvkbNn2d4Ag5rif3u0NUfjfxTptMUmJUBdAbWcNpIUvERd0qEmv49DBuY
F5lY/zKlWS3Uy+tTrNculGQy9gbUvXc9XSYAxh6C+PC4TrBJObyPrZqAYqWG7CAcxb3lJ9YNoqxR
hqmUidmOXD2CIgbJ0rJD1IJx/ZJ/Uh1Mtc6bh7sCeULR+kG2tZnbn/q0VoOvknCzsutKIBDsBW05
WfnnZes/GJFuWUWBfjBvx8h7KY23BFD5XoB1V/nzDDUI/2q7UvrIuHy6A0gAIJBvG1WOoJ8YFAqu
wAUfNICwNmfW86cmdBfpqw0omiqFYJMlYadEZp008/jFr/osQ9eOE85WJWziRa/DYZNprbp5D3EF
gUe7fidZDz/MfR96RZekLslN0PthnU98ulZkr/fsDLRHMdw4fBDGkT0fehL0HsgTxPCO4owm40NA
OupKd01LGUpjoQbdBZGeARc6wixlkFOQJtH2pAJAD6Z9/nk3kE3hrk55osao+5d/ovaAErKUUeUM
CKBlJTFfpEq6uKxXi69oG91oVmfZL+s1eNujDDsUs96m3kWZX3fL+GR1tO7Xp5iiyaOaY/jCnLc4
Is2XWnf/lXHnaopnhstZiRpHKCQ6NNxk/J9SbL2V22kheSPof8wfpDR/IhzaFcDhDN2fPujrSJTx
Je7c0kpAUdQRcwMQ9XSz8F5lkMn1q3SkcGjZCFO7/pBdhqgEGSzNaApCeUXb/mq2ovfatxKW3GXb
L1HacnwdjX8sl978V6k42Qlwb8kvvkOk772eEJGvyMG0vAaCzsR+4Ctzm4iOHX4QgkR6cuOSk70O
3/SQXaPgoi3GYkn8MmX/ANzLo2ESBX/NLTeAsEGjfTHWwMrNV9t7iNVX6eU7KUdNs0P9JX449Tu0
BvLu77iaD+CHB1+sCeQG3sLizZfsQs07wi9s5YMESGEnOku56d1orrqg60w5DkgRv7bSlQuxeRIq
+dVUIU2JDhMXB5gbFL0aJpVWcpxPOGNsSjAykIxA+eIRp6WXEThKehNuYOcstTLKp5f2JbwatzQo
hznaQ0NtEMH85ATKtbIqLeZ+IbvWt8RhPEb5KU01jwOXEQvJ9UcnG4Znqqw9DRdjuk8eJy8HdTYZ
Rcu7tGDr8j4idv1FBgSnC3NAAUCMf36VuDs+9igdt2pCbVzahBZo6j6HS2l1zaSNIpp7Uz94JBto
KB4kH4PkO3CsjvZ9b+/Sv0s8sxTI2GS63VqoY6gsT87igm7iH0Dc9tEHuHlwM43hwOJUtIwZjlHM
M8o5f/4VBoa+tXwkPVFJbkCfxbTi//aDCBrmood7lAesiAqf/QaDTao96LfMrjTQahkN0ZyM9xK3
kQpSiFxuo9rxpWaTeMl9QKZ6jWHBWdg00wR0XcsQbHSbuhxWlroYbGrA9XcQVxUcScQ2S+t1h03t
NYh789zmeO2ToI91tG0qMNGuE4y3vM7zg1P3ucKekR9I1Udoh/i2YQ3QAWvDg/6ysWUlvcMtCR8n
sCU9wic3GM57vnM9YWTjIMAzPGcs3f1GKESPlVq2MQd1d6ox2QDGWFSLdfP5N/2Bm0/5iMl/A1A0
kT8CyWp7/KLEA4CmBIf7WcFZkdu0SIsxZhGdw1BUEqyhrKm4DcyKDyancAfdqb/Tx6f3eMszV2+H
vF0KEnJJw7gHH3geSZZO9XvcQcPrKtrT9f8bhRp/10lEy5yFUSELpgoNQh1SgVjpwRUDHuOtQV7D
ETXHWLwJyD9EnBHSvv+kI9pTdSjClsT1tDxNox7EYQQ8Hrel1Y/RpA5MTC5LHYpI/ROg0E83dx7o
n1Q9ivSgIc6TezrdlgLRUYGz5nkxTvfkF3eEgGnI7/+CBBdZN50WocUOthEjatxhU6Dfn2QbjxP2
TzV0LIUrDcqjeZI2dqzpsjsx0S2Wsh7KvsfQpCkghOsmOtXNRxnpX2kxBlJl9pnnl/uzZuwtM1Yz
2St31vA8F5stYrQ3QWEWbowGyxLsnbhcQ3VjFDxnEWlvMha0Nw3WCyxkAEXqpNYHtl2A4Do29KE9
0gXBWMzx48VMymg3iSrUyP0yU+i/O3b3l8+de7mFXYvtjiX8Yf6yIuAnCzK2Z1RboQaJk7+pn9xh
cEolTKfD1zxJ+TFPfPkla+inVgKXIElyw6LKK33eUF0QI4bIWgtdpaBTTNvvNDsxo64VdufQRNvh
iMFwd/4p8MbwpsR3ZJLs2tu8fYPV57snftrq93eVXaGXbtwB+T2Z1aLCaLTCA8zYginzrU5ebzIM
Uhe8HjOQ6Hc2Gk80NfAb8kRoURiE0O7He3xHAPpqs8/mO5ykyfHjP8HBS7NURSbt3K5vRAmGu6nM
6a5SRJ4gYMPmp5rOAEXHg1Dybiac8VjkxoNFiLvCg3vf5YLDRSJgFDcyF/2uhzr0n+5q78cMLCjL
LY1qR1C8nqgrnPBEIUicRAoFQbEtZdixNF1ddK8RpQFhjsIQpt2v1GkrHIavz4/2sV1nb+ccvuxW
VRTRjYT6JN65zv3A7VTYKrSZ5PBLamvwNjSD9c0kysGPxOPalSUxb6SEOQT5VwSOCi7fm+k0rdtI
152aKJXuX9jHgPzaCvbv9g8Bs/Bb51i8Mz0oLDheigkN4JAt+QbmxACJswfvO0nSeQTcbMJMrtkS
/BVjN7KulF7AMqn9fiRbnhlQo71CQlnDMWPTDE9PD4yGFznxKgx6baSeU5GbjgA6JnVbTbnZ3FOM
xakVFkHOCShXcsTC6RU2WLNkoIldIX86yqlHFkNljqiQfECFKWQAjyJKVjuf0AI8N4v6/BdFjCfc
8ObUT5qHyGf0jydZ8iu9SwR9mz4S3LOJA1d24PHBvh2FwjzZq+w5gfQTuMrUBjRMROuG2bsIwX09
w7kl2QuS6/7Zx4/ER7U9sla1jtJxAcbN2laUDUsmf4awqJhm4517wARObl/wy46q7EFJzuS69cNi
bc64RNekctZXJmgfIKQtsr+cQtv05gamozk6jl6cPwzDzCMHwWpKJXKAbsdMEBeZQrO+lqPEqjG0
k1mRW23AHD8HtHTwOJUKjPacvAkgRohxf+zm2Grh4fCeSnVqe0x4VxTVdorhmC/Ti0Pivhri9U4i
BoLbybYDt4Y5qMHZGvVl+nrN81lWmvCN09ecgsRiR0gajv82fPec36p6Zm1fvFDl34hns6v++Ny5
7pFR775H+Eugnr3PvbujCz72vOVl9Z1AcLF/BRC8EWu6DqP9EyNvrCV4AJz9BwxZ4F8nfQ9SUDAu
lD1eJjcUMkiqhw+BoLUYdWImTK5pDEJ7lxDsEXszWvsdf0PHE5rHvse3xs7icG4FZyShYRBPE0hA
4V2UTtucCzMOynHkdu6Vn7RETok2FHqjWwTvIHwMaQTz8BolNjdumedRNndV9jU2ugXcCAUqdMIp
AcmLBZprDSc99MtxUpLjQON7qmnlDvcO6e48q104UJu27sO4R2ownnmzxfV12M3MmJMs/CJ+GaaF
aRQQdMIk+jlsrfp2OQ+BVqz7ReblKqBF5YPdcewsMlKVL/sq+JKmF7eh9l5MeaXqWPCu9gplaRDl
NxHGSq55ZJqRC40t1e14bYib2s36VXx63NsN19lCifyLGYCpfcDu4kLdFRvPCTj3rRhM4KSgl1rp
Q0wT/dsBIt9SWXLkECfzYoObs7HRfxQI4s6Yt0nfFffRH+qjf4qgsI9o8s2DnzdhQQu33C4a6pTO
Ue6Y4+iHU/sNRJpgDuXogfoyE+wXgsW/odwM5xaKZ0SoB7ztjQ5DG4zVse/oC1ZynbpTZS6EG1hD
8syO1G6dk5J72iSF5dJLzzC8zuABi1iudzrJSVmfnO+qc5MX6StJDpqzLGMcOI5ctECP2nJt3fw7
6l96SRulspyp3V9rZBQC+tpMPOl8EZ1y/kt0RlpoVJlXolZbtpeSPRSmQxLFqCsYe6NUERsYtdTK
SQ4cE3NzcIlxEzYoDQxSAQar1N33Mq1LOgU2byhdxzyERNZYRz+SSzdrw8y0rNJ9h1or2/RVntti
MCJxJweK35m6QTE/UcENf4AGQK9lkvovcdktVVfThLk6VesGYoaP/dGSQRO/RHKTvGqBkKPDY1E5
iiNYKjcA+4rj/nk2NrVBDMugrJkhAXK3PRzBS3KgPe37TzHvd1xVyMdllwroskwWqyiqDABz7dPi
rvi5JjS4Vspdx1HEiOgFGrYCxzipxcVYWvGBh1GRP+Y0vNq8X7nLeK9insp4NiiKfhGtjr6mzKe9
AO9B7lSQFkI2owZHAtnUOnMXh4McgQEi7zPAVkN/ZI+xrULBRakWbtoOV8g/Sc16d/wyJZstjZkv
I6qVs2jeIWwEHS4bXau6+YYJ+zsy5FrQoX5k+69FIwKkK+d0KY12pIRtYcYGj9h1+4j9RJam5rMm
7iTYv4gPVRsHjc8FrMCqwwJwGamXxxDI8mEi0SzwE+jCgKHksPpMBMEUeyvcIuyxeV+IrTnI/Ohl
20Empr3+Ajj/UNivVJ3G97TqXS7kC30mJQHnwt/4dE3pEa+x2UaP82CGX9eWpLAkZuMUdsPzghaN
ErgGnvOHKqLATgpfQtZwjFKa2XUGISw6EBA+xz3yF8g79a1a1hE10agTKqUkgm/wGBVyItKQrQNB
3DbusExfzz4WXVN3IX3HWNmuBrsaoPVaYkjjRJjO9xyMZRzUhEuCJHH+j3uy6OvwqclQCghR01BP
Qrb7ym6xliwJMHI8FqynZu0S9RJU3pV62EzSfO4/+dmdHQMC+iyZs15YOirz5yY+5/iXuSvs82n2
W4VBDDpCeTUnm7shUcr5uK+O1H20SaHVCeC2GsKFt/1eUItFICYi/CMbNBbcv0CcAUqbfOyz+vFI
7VzGHv55kM47cvdvXqt4j236SIitBDmRfXNQN4cwt2kmmcCUGrKNc8KJPFsb2hWZSPGB3YcXlmY1
YPwUIfjMPJ/YiISxH3jXHlBP1XiKMktr24mul+I/6TtUOJ9fKCDtRrxr2quNU5V53gd3oMg/BAOm
KtqkeX2DNzRKGWGiMc/nZlak9U1yEnHUH1c0PwPRUaCm1CZ4HRD9V6cPxtUi4cIEGkdXKV8jJd9L
aJkDkdl2mqQ0Snw2Z2Whqc/V8TD2Qg4JHBCgU4wL4M0/zYbZkAviVZyKxYxkZh2Y48Bzcz8uTsWV
WoMWhlaqxQOzSp53MKbc+aygsdFHnetO8rlW3uzsl91rwIFccsD13l/9DtGZi8kC0bm5tqY8gLG/
4LGcsoUm6eV0zYALHaRbf1YDH03yonjIZdcdqt//ss3/3/NbZV8mN+jI+FHPJtWho572L+RMkq82
NYQ8nc5hwnSIJ1LgtsMICM3ET92jC89+OgBQy9zqbYcFVbDWK4RxL0fNET4UinxuT608xUxBO9tD
IdhAUepptqtyr1bV6M3FAHsRRfIeo2mF1h6iDB2FoQcBXC8bP7T7bG5cM0HYepDuq/lNbnd9YDYj
kRjvIkBhc+74jXtACV/DwzzLNEV4G2no7Mu6kyf8C0Sv0QzcRABYp5Rwf4l35fUwjvr1JUvQDHjZ
x4+SWilFTtDtBst58pAI4HYdv//xpQGFT3H0ZB8xTTCP5/qGSbwKV40+9afMgmKuaQcYQe9ySp/E
9OJTm3YIK6RN2L7EAYmDfV8kg8GAEXnSMsTB23raCclWIwVuidH682tuN0Gg3UYLRRrUqGWQsUiU
5xGouLQR26y5YNDaVrK5Ps6OHp/X5Y8XbOGqMsXpnK+L1X2wsLyb8KwiKopaX8W3gIWmMFVM3hsI
Xj/DqwL/q4W+zWyJm817j0BDj9nKMwsG85R0pLL/O6fg+zAxrQM1E7c1MCV1KBoGJueYBJJ1ny8a
BV9o2NsqkMoThbjsCPTWBO4LUMyGrc2ZI1EAmHsp05INuyC5e3LmR6nNqL7x229ndoX4i6UcWGkq
dsuWtec+aWSkfkPxy5sy3AOShkh8BZlEOQwbdyIKatA+KjwLe9yifvwpyh6EhMG9wWV8bqQextJs
+VBl3ClvVk/ZLPRznyjzJpqCBtia0ES/P4JiCfIt6ok6YrAZPzc5pIgZLudnPfBWJKFgYw5oihLI
uPOpGGJOF6b1KxBKBCeL6tnP6buZRTd+ZCiEOtZhUUyuQcBz550/Wmo3WNC8sewu5QV7ecuqd4vg
gjumU7e530HKc7XBhQV+HVlnXcsHg+iFydmZlJtWgM0anzGYBTmdYQQjezAP4p33V0KiHQGImByN
Q/cHaajuOrTzEr+vYQDzLVu7IZMWzzOrMyPkWkw1POkiH/axDssZCqRjxxaphVmME3cHaZmlzJty
jq6AFPHJ0xyucVI737hFdfclvdwaBfEi1AlK2Nmh+a15AMQtvdgciNuSjy3bvTDZaXg46NWN3klu
2414COVQ9sV650uqo4BDiaMbYm9LgNn+oca1MwerK+0OstnTKE33Wj5oG123lkq5Q6RgxaDg2Lc/
npI2Gu0zjUvrdquy4W+I6kpiCxJD/Qa0xLJG8OByoU8rThjND1yVEspFVzxsXHwGGfybhYe31qDB
iy7uzn2HFFYK2hBfs7APpHSO6JW7bBmxAr/p7OuXQeL2aznVvnfjfAZ/uVgbwV2telItkbb4f947
2VrVaFi+HtkJnAfLJc1wJF/Bl9yKnNe1ssKbcGFYl/TK3wSrifwOLQRfj++BFFSXX0sCi2Kuz158
qkNhDKGb73ttfLKZEmW7bLTbtLZ/PS9cjtcNZaQOCAL9pgeMZjebiWiUu1B5x519KpItHYTqwp4S
okByumbvXWKDgVOQ1SZQVI/IVHg2iJhgSZsCTrkFV2uWY8j/TX0wA6B+3aM0tQikaGPduPAaA/sS
B6HQ2HJoVZ7WHXxQIwrQ8y5pT1kntg1Cnl+A5qPv8iF8WgQuLbc0qu3FtUJB06kYFXgvXlme0hvn
lfWZ4pSfHmleRissoIHTvq4Ttqbu8Wyc2aHaAF1Rc10p0gc6GSxtPTYv4eHakvMBgN7W6F8apIyz
ykg1yCzTs9/KPFYkQGQPJKzpGgt6R9+ztPPzby5zwrog5vdcpDtGc7Pt1dN0SXXtkqEtpCxgp6Hz
Xbtrqv4pMdDm8M4AHMKMIYoQBf2huxahqbmkb68Y6/kn/IwsUy6bkn/1jAH9APIWXbIOj/0jd2Lv
u1fFT7b83ntnLyf8vHqr2gFTJRe7I/h1Fk42XAVkZiu3QWwPERmYFQr3gWx3jq7nc76WpFH22OFl
De1CF/Zqo7c1LrbJXeOZMsalskqdxEciLm/QTpoYed6Zf/BZWR/prjGgs+AZUhpiJny5rW+htooh
mnT6kOiOFbI/MRlFC9ejpM9CR8wFh3uMqS45DMA72hHCZ70CbKyr/QcsJ+8wyU3G3EvBTEWFxfNc
ffyYhFDzrRNlu1VkPMbwErn3hMuqggj1gs3kWVBB+CYhx2OxwE78fXgWf7K3Li/Ru7d1iqa0XN3b
y7abohpSP3Ll0O03EcrTKqCzQtRZYPLN4hMUMOYKf0bwK6qBol/acWRFYAerqCFDXtDi/F5ydN73
6gSZ2Mu3KE0of05En7e8MTH+PkfE2vEIM+NYPnvJPC40Ctq8PpVxkaOEF6w2OeCpoq/3nh7CsXfq
YPGt36SderKnH0YdFaBxlpXM6HnO3Bt/I31lghKpFwP44Y4TpvLFgrWcEw1vb+Y1u7LawBCBV8do
qE3S1tn7cDyrpVLSaAvmNXKRRSjN4sJknsY3ONYi56s5AO4pqq+KzWnNS46SAUnTYKdX9f1SYk0w
caUvs9y5FRMMMIYWOQhcgH2NjCKqbp6s7z6FS63YSlV3ZeY5uChokU3zTtBMiWzwej6Mh8m6pgVs
NCRUdpOxBHvr5KNPZxzbe6wdKYXjmLxvgGs0zZmFHBFbVlOKLSbvvzLcGlFhfa0wAeBCv7BUmhCA
6POlp5tJClWEsqZ6vyJakON0lIkWJ8zcTex4lMr6HNbaBy6FlttkvlInJsggPkEqYIub+tRtwubx
JpoS2nPSR+7R1qEjETBoHj9fAGkTXjcgDkUnFsN4mYx+OW4O0FGu1tuYRitCw6XNiB23EFysz6AC
urJpTAVF8UpYAbnWr7faqJi1+g/3mDgf+sJmfK8PrPLUpt5cc6+6zBHHIWFwdIE1MvcSN24Ru676
bSGtaY3ARtKemEo4vWF5CnU2XVafzJZsQ3B6QJdS9bSBwGuONxl70GjJDIPLHxQIgln8I8Fz82dY
V/wgGEV0qiLB+mMEYdzsfYpcNLIzPKR+siMNc8Gb5z+pXU3UNIwhVYf089OIASk56Tq5975lCoxd
WZbteyQc/m8l7bKRbMg1FXez7Nc+qFSUTiJbAs4cgl44v+UBOdtfGTf4zWKDFmGphtTrrFiv0+0G
gDIryoMMEzJlv/my/i1/frtmTi8rfAGQijIOlK/vc+msLeZoouYXjvB/tVWM8bCwlDkG2nj0r5D3
/iC74NbOallYCf3MzW3zjgwLmIeZzeq/p7jUTR/OalZk/5ls3zagG8xFOqlC8glFjdfpIyrBwlHV
iFQYKGnmam2pdumDLZu5j4iJ3SaHpLkQ73EeQi5dL4zn80y2sf1BKijdH78KCQBTUqyEKJTdjwgZ
fQO8wBPBiySrDcKKxK3Ihp4eqr6SGIhblPqUqL/GagZB8p/AkGqo0G5B7BO93HkPAf6SKwtSOA+M
/3MJfRXxdHskwpzrk0vt3gEonm/eP0GTntW4guu4FSdd5WVegbuR9tqxBkACDYCnUNKX44XdspNz
7MJ8+oA2M33wa+G/EXBU8VIqLdyUujeZ+oqv75ZRIeza+sJnJ200pNq900+DaN5cClOZqAAQoJpX
LckDsFmCTLuyqHlx9uH4/qm3iY9WUOlQgtHqpvwPZMEzHlQTEJC8ZAAQMYFeTrdUoy5YThex+UwF
oNYnyu3IDqdGal0QfoTZ7pKVIFkETfy//WBwc7tySr0yB/X3Yv6V2woNtCUeAsMN920Li4FmOXYP
zHM7nNABzdeNgtj66M7a+tap1NMrTelPfAlv0kf1c3JGHXUX7mmj8yev8FMgrwCP0rJH9RjTtrLH
B0mz/4K5mCV6nFAFgvgkLRRjVV+q7kzXAfT20vt7lHUKEqFqbfc1VVI9E5kCgg9Kl/bFO346iT/N
WYHHs9Yt31fmy355a1U1iAkESyruPFBnS2dh61SsjZnGeW1wHXkKfhlaH10EVLIwZ7jeJ5GK/uBd
bwgeEawxkJ5GAHhNHlcCnnkELd+jftQCYo3EtTFBnlysNX1ZcibhNyEh5mOJmzisDtrffLEv31xw
0AsCI93Y+c8ssLzy4ssNftCxpmxVOihvWW1mUaYqKke/3si8ADOmzP6U0PYrKkSUX87KYrKtwDzU
iPq/rIRdeghVWJ4bU5hxylIZFWW/nl/cyhkCKnK7ryH3WMwRpPWOgBitEfd9/tpouvSMIS1CLCku
6D5nGVr9ssYsc8I3/v/OMbVJ7qLRnyTOSDfHGHf1iSr229DA9JuHGsq85JMIX9QIfHSwRq7IeNo5
7KT42Tnuv+wWIJgtPHaWDRTiimiTIDZgyQ3jC9SMOmC6/0FhxvOh0nrRGcEKqItnVK/r16YHZPkk
H/KriHz+OEEB3FEDJ3LkjyiDaEy0Ad1PooS1870y4k6f00zoAu79dFknd2mYW/eBogwuw2z/051l
belgIyj0u3YKbPX2ZKQSEcCmFhEO/OAf4T4FzAT5EdWM73kPsMzl1xHEpr15jUiHw9XoowDgF8VC
ynDVHraCyNrDYyUdmOcI94Ra2ikYVupZfQ75fO2sfOs2Gwe4ZX5FQfWa6wTo/DHYywI46r9wnEE3
QIxcErdSlMAsOJ0FB2XKtCpbmp2wQwj3zN2Qi8WU+c5jdukqlL/gxnsYLkZ7nf3bi5o5xNT/3wO1
epqKTolmVXDXEWzHub+qfd2WpZSZgTQ6b/XGk5jm6oJfX1njg3iYD8+9+dOya/YPl2t4QMaZmiJe
+OGDwhtmVC2rjpJlFrD5qTcxGNJfD5x36tkymNY+uLS7TcgBT3VSjDzKOH6LQ4W77R/woF5yu1jE
w+w16Lh+PPG3r9CsGIFM3l7qR36pJisLeEOaAHB9kwEdKYbcSsHxpxROZs+zNJBnESDwAdqVPKfI
699PGf8JMpMAIxVreWp/yA+zueO1ApftuLry8rAS7AqYC12Wtk1KWZ2L5ZnB7uQjhfYm+7QqPqcs
L9+XfMzbfk1Gz0HtPZkMtDyCwOIGszHrmu5Yyuu7zdf4D33k3QTqCyGRLcq+nyiCOD1ss+qhO3m/
+47XVWirBxQUb9wNZhyisynACXs2kTpE5Lh1e+eOXb0jKHPinGOzt4eovtQCJy02hXA7HLf0/p90
irr01d8ieYJq+9EU8qG/l8Ottenj+wIDhSPc83msaalbCEIZHYmPjI+mRUJefoQcf3xwZviQ1pBv
/u+Uj2WONdh1jZhyRACKdOaX5P51L7JSVuoX1g9/GXxgC24XSnrffCEX6s5y4lHbPt5BCpCyg0x3
1QrNUj+DfrjLgjyqkWKlG14dHmEXigC0jDmGdxZNrDUKTtXgt1YDKE7JOj7f6FG5+rVBsNhiHc/+
9jwMhRfb5PhOMvFymtvXcXIWii3BQJ8ChpAjXaKXfiSnF+gF5cvZjgpZlXO6qRt7x91mH0VKPcSe
3g9WlzjXA5me0AeICHOP5lADQyh0tyYPeFYP7DF2EmENp+sIG8DIeBor6rEhgwMzFA2VKTII1/he
xCaXD1VTi9kNSTv0jah4jVNbmWQnEeBw76ZwlQqtQI6bmArp86PCNczj4nQiSTcmLX/8/bbbwRc2
NdNUsj+anUrxoOJJH6OJtYrZr5RY8Aw6wpPyoAX9mieLtBQ0X4o0T+TKMe+wZh5T//DMKaSg+tfe
Szs7OO72Wfr07z8hq+yJwx4NsMNeg4dRNgkvbXZ6rdNsR20V3i2R+Mdi0m/+Lib2PMlzvMf7cCNC
DrF5NXaJvHoiyYBhApLbgqzaN/Hp7/vkL3TVFpt4EgwN02Uan1mCGE7Y2fkKsy9iv4Q7ptpYn1Ut
jEFyTb3E9O1w4ro/gf5aS7ZhU+0fFzItQwgAf4EZO05cLFs4vwIyjx9LHqqEb3EaaEWbrVhNswm4
KcNNRGgEeGWd0BHKoLpWPEQ3XuGoSyQTgtMzJmyh+e4LYYkST2pfzqS93GStRygFirqZ9t2nenCh
m0Jl5n8Tohv0mD6N42TrTJMMXVAYmWmAvvZnA7+unjocD87cjyxhEAWzhFAgw0BGLzb7MCAwE7PJ
kejC5TfHtQ+9JKtffXtqjk1ArdtiqWx415Bh47L5OKpZFegSuAXOqZCfXi74V41VwnQ8JP+DLi9w
NLijQ3nMAfhQ1PkmOgkctyQmNTCUhh8uHsMBVm7+fv83sFPPqsaUwgWsJXELihYGKbl4Aat9e7SN
NKwvybFIj1TmmHtE+UAjgV72q5RSgF/OIRVHR6LXw427VLIaMjM22d6SUEsqqZVUh4Sv0nEBEjPQ
/Y/hDXBLypPGSGSskDu101kflQpjqTncTchT3yTYz3CZOm613Ut8n0WHPPGr6NYuMSByBPpHtywk
PNALY6y+GJQyYAq/CowcEXONiyi1FNa1oH9tQetshmRNWZHg8OKO6sh+sfOu06Dz7bWlIAa/vlql
zx5uXj6u/heBsVwVSfeNDflogrBRCdtFvBvnpDR65pmOQvACCa/86095TryWC5XynCpEKDekUqbe
2FN24ADyWrA8VuICoyWFc2HFJNWVCXSOwFSahPz9Vd91U4q9fFDKfnJZF36TSoqFeu7IxyFMHXE4
UkN0uoiYjJwqHuyRe+ecHl7qbjTFns+N/dVsEvvaahYbNzDEMcCEFWSUgEslygh6H9qwV/24jfXT
6D/mVvJwNiuK0cRABkpjHF7xgCE/HmnywqgGV9+OOE+M/z+vfUFA0PuGZp3wOZT/FBwLCsg6ZQCn
9v82g9f6Nzsv/d1ewI5jbL4fE7bmIRZ8G7FIF+9TV0UGYeLpMbJ1c4Mdxh+yKHkt7UlHBTlRIgzm
WWgnB05B/Exd4ydGB+hVgYxnNNPcRxS0qHlVqvZDGNOoBhwzLuXn9cyx30sfWvCpjG8mmd/kpdmE
ppwBWGTz6OWkQi1zuBV25tvMW7OPJq7mSMsJJ6IOCFGYx8i8IaLA+HKwEH59syQ/2I6oXTQTSLvz
SxhAQt/Gy67Wu/V5OogQUQkuas82dsw00cfC0eOvzKKwGyz6haBjJ+HQoOQHQ3wWrGxOQ6npc3Fe
Wg06dHZcpyZjz7CDQcDm1kTZBSVCw9nP0+A0r90JvOH53jai5zqsTODFVHzkAcgd7HmD4CFWxsMm
NQd69WfIJEnhhmwOD5GLJhy9ytW4FTKNJacaKsUk9DxGwMbj3gLcl9YRVYg2daUUcZQ69Ax7ngtl
OzelR6hrEMMHK35WRDVxhosUTtK8EA8lOkg1CTGrHjiWdBN1tXiRzjYlZ2N2mzhs9LWJVacB/9vd
RBL8G3JaW//W0i6K71HXUExEpsW6wBMXCoOOs+s8gDm3bs7rk+5AKbrEghxydBrKJAH7XYkN2+kr
loGWwn+3FfzYBTt5X+l58SzR10oA42bqHixPqZ786dAQT2cep7jtXBQbYF6NIVe9ovAQfWNrJQJF
Lt336OfkrbBX3Jk3q3MAyarIu2tORCn6mLkMRPmR+SBnVEUkWkVIlgQouVF7Xl7Gmh3761nV7PAy
HJ2GZhR7mP+9pX+NdGAD+CuZb6AVX7FmEowS/Z8B/cmsxh3/e5ei37TuYlI2AOPRhgqgDsYgTa02
ABlwgFwceuVF85Pk6pIggnFZ0U7CVCyZDEI2e36c0X7pVknf3URPloFwiMRbH+hgGQEPYLXBqUDX
SGdf444D0x6wiNPFjIYosvN1jPgMJOfSaYryke2lk5j4al9WNItXhGNJoSPkJjtN4lai7FDmdcmE
oVzRzsE0VkzGEsVgeYJO2j8Az1xpdIKKLDhQN9xILblZLFD1jSxiQcIAqS4FkdI4M1KXrNLhZpy9
zCdKVNveawU8GLD61OYye3PT+Q/s8lp8RSar8AZxqLotiM3GuK8WGh1L4q3F7vUIMYygVHlfpAaX
PTWqfVDdT5bjZklURYdWSsrs3OvjC1rEx86HX9WCfhWn19QjUa3P5pMu9E1RWnBRxNB7vW4Z6Hef
ltCz9nlX6f1Yqly+eoHnxDd+n923joxk1wuCkuhaogu0FGzHigSGCJL8GSc5tcXarQdmiyU4+GFT
nnUQnvGZqExrnoL6+UpK8WNGBFFntqNIUa4lF0yDHa0tdIZ68mQkk3uHENCZcgGQWnn4ERQLrC8x
JHRfAgBxA2OnxvUUk/EWKqGY9xGlUicS3QE/PJM99uuSTDg31miyg9p+590RUXiU8bH78Lha2zpJ
vO8jHHXNU/A1WRQCdh/Ke35mS4fuu/d2wipv2x2s+RjisWP5CbcVYR7RIObfQQNee4pZPD8xcMtX
d/x3saddSX1Ej6YDcVXTm18D/laMwuxbT4nWlA32g1FJSB51yM+gZnxbNuf/xKIrxEHhfaKlbE/G
PrBe+oT4m5r4OqvN+07hOj0Sfk9/4pd81BpC2uAvfulde7vdQ5yWjMeo9uREkRlgkhrDf/jE/+8J
giqyER0j3WnZVylAKs25AbwDYP9VcrXBsK0JeoVYGGbwmhtX6SNIXadHFZN/wfDk9OuzKAEI9X6D
iiz6bqTRtq2C6YfmVNfMyal6hUxlA+BIEk0klhnzld1REOHhr13o+PkueVviimCq4Dl1ZciK8PUc
znqUAPO7MbONsLdPbYtotuiim2P8tWAX7GO4HXg2bGrUXLfabMXP7tWdonNk5BIgRC2ZejYPWw2L
e8DfGRGqFHZ1r1VrIoZd2MGbx8aakQnfWNuPULiq4qersOIP4Ucs5owKTycnhG1J6vGkpZAG3wg8
OYQH8LlVQQNZniv48DSzhJ1pFfpWUiRj5HxsUkX/rqEkJXIl+PTyerKsfBSGVGjoGH5KX56F+GkW
sEMSthkpWNIUW6YlXdBuwZq7Uvzf1ULj/sQTHPGvrunoAUl3gRq1FQ566CBsOAvEdntnGeggFY4q
39l/N1c2wJcd9v8obI9xIAHyfJyILqg0l/2bE9CSQosok77A134IMOudd7RnjdC7yh4ZxV2dsvF0
h0Hv3UF6URol8UFUFiKUjAEzlYw6fg0LGRPHJIsDknhm1L9yqt34wxk0Knky5moOkCJhuiM8RpvQ
M19gk6MO+zv5TT1Iib9904oEI9Ww3NgfvYkC1hTfKsklNHRjWtXYJAXxlWSGAolslmbTkGyRbIqY
kWJVhaw7Nzgjy16kVL7AHeLN1sfUVtvyPy0hHw+jJjyIbo7uaXgpkqt4ZV6dfYlDg6Sm7xST+Z8y
tG/TiSJ/C6wPlY2CqrJhuKdI8+iENbY/vc6jW5E1v33aCjX2zdUBowJs/Gt372CBJjzZqjdo4rkK
HsBKnLobkn8SITbrcKjW9HLjvC+46X5WPotgzKNdB8T4AdeIwJrIwjNuVoKeyL4B8IgphLrZWlFG
eF+QAqWfjY0s558mjCvJZivnm1bDXVeTLcTUVKGvd5L2nGlLTMe+fIIbq+XoAlG26EOeM12QQhqP
xTmi6zwGDebV2V9NiAQ4vjdQGwwsckedinHgGF0I+juovmgTB6ZINdb5dOIXHMywAT8gm6aR5gYl
fKUZ0dqtyzj8S13JbVpLicn67/q+2K70PUSOZkK6cZFRt8MMdH8yKGpo01U+jo89AMpkOjtCHyBB
GxZgHnmPK4Us1nCtddNzNgkyhnlK9RPUkRf/sQAfX9xPnvyvJ93JIBYdyh7rBMMWCbl02z97J3O/
rwsQ6gEhMTUikagnTM5CMq1GwTjyInW0WbMQyaxI1wQLobtWyKVoxtY7+kQfYvlKIBi+QUKtcih1
ut7DMx6h1WkEF7X/CDwBI0kxwuAMzGJU6UA6L7c9Vg/PSx3eidfeo7Buz18OxFIBezxeC2frc4+8
2reqFkboLuq8rNmAYyYFbCSzo7YQo5XUY2hdaBzPl7+6B/4g2FDcy2WOVYy1NFxVs67KLRMUDeIh
yyhMeEvHASs9PVw9Si+HaIHlJ9DKNRySqBB+3E5n9ZGEYMqhsp7JbkBleavMEPDaiRTMf2mmJmhJ
VvByi2U3lUEjOQF3T13vaQAnBUy7Dl/dOXhDnPNr/vvS4fpLvKfQoWMi8S7yGKWSUC+L5RqZs2Rc
cf5/Zs3MlTMcIBoYCFH4zNEBjc6MhjaRMS/Qw0Am3Yz25HaH4IR9K4/DjJgijt4zU2iV8oeCpdCr
oChHGGcKo7s29/nWDbRKvlfstaTveOQW3jVDYWDMRPS/tGjqP7+3fMcSOVQhPx2XMc6w2xZJDsYo
pORFcy01q3jQsMA1WH/ZYSmxNcVvYwhFtv6aZKMgP08fgFcK/z0m0196XNoXrvffOhJFkW8zz5sr
mqlUoi3OUyQVcywxckCGCx8vKlzaySgUredVV+GJoaarK7ENlfOzh8h2Kb99+cGPSZr+nSVrRl9p
3bXqTCwYUTsQIUmOzxfVImWhuzIv7HYcRiTrOXDy7FtPIO3a9p+zn5zcrpDjiSJRPuPorFKNeGg1
nu2WIkLl1J8P5jHSASwp5phavzrhmP0gGkX59rgw736ImA6JG1z6jUNXp0dt2EmePPTztD4HiAm/
TgP5Dhw3uFwKuC578swoRmWO9wQtLw8/db1IVGeIKcJNxPu4sr1AJs/Kx7RZMgZcoKuDL+UnL04Q
caToLPzxZXqTZm+TpF71n8MDfUKIae3/wVN3Nf36a0TXtZ5IpXzixcNIjQKhEUfYDfNUrCTsipnn
5LzLPFcelvLWDI8xS/2wTLZ3zOzi4Y9tLabFQ0GXrJnQUCFG4MsqrcRrmbMWVqwP1sr2xMVqY4z2
fcLif/95oNQeOzjmNquVsx9nuv9pIYCGhZi8c6db80lATY0pyN3d39g8A0sk2IEoVY2n+EjSKS9U
taO5aDoRRgn/6U0fkoLl47GdQBfeyQdnL6PewzmCU3fjWrrfRgfIYzDTjXr1aB9Oyr5a+F/4pJHs
r7EvpabHlM6BjS/B9O5IhLYFsyv442KSQVp6EiPifJBOxnh/JE/yCzqewJbit7hjJCW1i2qkHrK7
bpFRwlhaeBBS0J1/tpXU1GF+A76fpuOoZhC9DWT0YQj3NZjWD14kM2XDtQvDxapgm0C6O7nsfZ8s
RRunoNYoRdsqlAMTckhbAifJInbvQALb8ZtbbPH/r88i84OpAdum5mOf2oxEc5qYU5ArKKoYOT6X
epTvt6lonvJAmp+zgwLgcCX+VpKGeucYQkattpGUnI2T0p8tZ/Sb0NrdTT1/fv+nnwKb7tP7mEz6
YHcgjpphjvPlmTHdqWlpmBBSoS9dc+aBIbwFjvbTeaqGgRoaw2PDBAxXQX25Vw8hB84+onsL/cUc
aum0J5ymBMFM99KRWqBLsge1yQ/4oNWyycHMd50vGG7RKwqoWboFg06rMEusQTVb3NDYJCy5aAsq
QJg7VpADQt7n6q2JPBwCLEnUxXF/7Ef+rRVxUe5622Fz85ZRl9hpsQRshHLkMv22YH1EPu7p78LV
osqXMT6Yz6YyIPTsj1yoBpQ5aBeMfmUnpf8cFDaE7JAwMk+CbfxTKpCUEyD+ViCDalEqiCxOk/CH
1T2bhZcLBK6G2pBf+47si0tkUZLegvw04NrnMSJqV/j1CVGS1xzNfOI120tWxtuIQN/n5501HQLE
bp18XcN7QjLtsenTwbUv5Pxv9XgDd7FWgbNG7xxI0DDAx9TcXQkjEt3oUcgM0Ong9Sncvy00VfbT
bku0OYnauJrmf21GFKybHd63YV4EBaG5QRtGKhAKJgwHhme7B0rIxXv+W99XdDO9PPOUsmrdNMdg
5rufABrbzJ2RYETfVi0/jNEnh2vCaKYw6WbZG8EvgDLv3tHXEyu+VUo48cptmDJw292EU2tqy/jG
W+sUBDsb5YUY9WO/tk/mxwmX8PFywNoriaoEn0RPRXsNC7j7TEKOxpniAkWkT2jucJWApE4u5j1K
xXZ4WFow/piX0e9ZOltcjoQaXk5FoivQ8Mfr9mVivp8b7L9XC0UjkKF+oH943ordRIn3tg9a+XnV
4/UhXnC+kdUsel7CaunSZ/SKbh8xLksBjuPNe+/IzUHfY5ti60E37jfKjY+OlRJ4SH5zHEM4cUzM
rsoZwjvwYks/P3Qu1+Dbj4tLBLuIDpJZNFbDt7irCrjr+qEtuoXAnYR/sjzUnPvDLC82oBfDaj4B
+jkgf2kYkH5Y+6lx++b/qEFXDvdOKMD5opWM5zhpFyBsC+I6lc1p7Zon0ULIk0u31VDsYub2ioO4
t2v1Hd7MHNnTi8F3sLSGoSxr5YhlNrPF9/ecCTwFAetUJgr5fBVCTKDt8yXrfGK2MUn1YhJbLJQg
JTwcll8+2/UCXy5KdTm84OWF2YtEQxeV88FPmUnaJ0IA5/ggJcBwhJb0RU7IOyUeMVFGhcRyUV1p
oNItVp8AxtxvDp/+FjUYi8MWnx7A+yjk/T0PLsPVrtb477EnQufQS4LVBNPflkCxz3YzY+Ic/XVY
7CswNiUoh11ig/2ULpmX99BKMrsoEXlClq6gsU+Rhbo3IxT46JhVytS73wlGzxKhvYDNTQlxTQqh
pDDa2KuO9g6S5xebFd6+kMd4NVnyD3kx/nmNVio3jygCg9pD6ley5P+nnak4ZShrkgxSWZ6+B0Nd
W3aeDIUKQU5wbMWzKo1oQ8/o869FShE93ACd9HgkfURZW8EHNYESck47TSn3XbEXHqPvLUnBXgXp
69Dcu9ubbbEt4BPWIE/lWnS84gegSu1ezhEgXqp52nLAn1PoOPwHicAsrcIqfXR7yazV4vZ9gL4U
WzLEa2TvOPZIHOMKXSUUN+tFfV+5qMlBDfp9k7xD0pwfo+FAjNJHy1Ap+IdmyT9LYPf5tvTJjsub
jMx4EiIFRAomV2rxlU3BjF1QC7UbbDEwhSXFU60vV/VsMMZJEsx9XPE0MCWSjFQLAqhx/CB128ah
uXbAl6va5b3SkTzXmvSehpx1ApCMiwHz43d2R8CPEjHGEfWx153qk2fwKDZRp85tndm9xPDldq6t
TzyvVw/HnWfHWlgaxyRh0uBY3SPQBMGAETHSXEFq4qR6tqd/0huLfo4STDFkXgvzq7sszITiWrj+
RA8eWg/iCn0mczTWQO7c/aXROZ6cJbHn/Oi9AYqtnVMboBLrFmYZ0i+RmUBIF9RqvfuC3JPdh+W0
hilUk0KGMzn5wEPgbbE1cuOpk8N0R2nmZ3OK5W0h5eAikprBmZHqHtnRhb21LpF1rA58fGZz9Eyw
/oB0HNRuC3iQM9ndaiQwoxH1wqhdicxtzPBLvDX6BcBliIWufsu/1nTDAfhyaxFulmws6st/6uNK
XhoL4C+N2yxBp3AxKUzeJgeed7NJD69tbhJVwmmaQgaroRfUv4U9eI82Sf6t6Q/ZloGSlNVwUyEh
OCS5X5C71MRNrkVwFG+4aSU5AUHDpbVi4m1dnaIF0/RVu3lQ6FON87sGkeWc7Ie/12zGBa31EnH/
BqOOmdhXmVFA4Q3aP0kIB2E8mPLBHanyHT1lWtEWr3q18rCX6VEo7v8b11Oa4MZpA5BzKpCNYBGa
ViM70lUTxlkv/NcXC+bHEbhelca6ijKoQNz0aO7wWMt/c0zW21g6AmPf/V2AadIpUM0+rqEGX0cB
jbu81hwdhP276JCOJcFzMwbOJ2yGL47rH2mJVxIQDsGfatWm9rVYwpjQuJ7yVtuJT04ztCs+zdA6
DVzvyYwS6SabkRhaXiTYWr0MyDSCIsl5TIljhL+ZpEPaofJzDSOCHwhw7UuBR1LL4YxEUWfz2C4e
8sEkS67ZPLFC0ProUVmkff63qI41PQXpnb+h7Q+culSZgUMV/3pw4khkzYtKYI3QDSHKmejuNxxx
XDOFaPw/LAkGcIBTjg+LTVzRfbFIMOdY0AWJj2x9Dv+w70iCnptIWTdI9Uo+0p8wvoeh7zCKxJB4
TGohKfg4LCnK3kx8c4XbsWhgiXvUEDNhpWm7CE/Uqx5fDqH8Nr/RUk0RLIJ55W1YJN1kgEPu4gn9
jsQtM8qpKzy/epAwODvcmniWvWfruldWA3JuGLmmrOPeu51GtqYGOZnKTN+bbbPeQrZACfILB+9S
W/RVafuvLpsncgXQRKaO3Aooy8kAe/sL7UB2XhGD6s/Y5Rvom4zfRlnz3nHjDuKHk7bDZIj7OFLT
fiZwWUHwIt7xnL7DxtifzpQnJctbC0+Oeds1caSdSJwnjY/PxYRDLnNp4qIOr30y+6Uuq5TQCYIj
eS95UsU6hl2/i/4pDjXSizR5LRM/waGnAZzYjs+rGJlIoW1Ks40/LlS9epEOVdaKmhS4qre9yG1N
cVkR0CW/BvwUwfinTNezH+XVzu5LT5GuPcqu6zshoGpQwbkhw1JyH7Dvo/6CSpiXyyyy9zaXvbhY
3UhzJHhGOgu6LPcxXrUXU3CmpqfrlfNksuI0zc8eFWOy6/2LD3Hst3ldt+sUbEKH0CDOTKuBHDie
O4ZPp3C8S9iUxAdcteV12kq0xwY/RonZ5KeocpYxk+EgfEiF9tCpb/WQXu26xarFmSxPaKAfTLm6
0jMwxlK7yVvcB1aPf4D7BUuPb6dgKjNPa/H2nFpmrZauxR2dnY2eiwUzmOYHMGBgwY0nVIcrPs2X
njVegRdTNiDmvd0qIMwomDB3s+G7vxVPZ+QenVWT4jE0+eQ7X/Gs9yXv1gIRh93SA5T2iQImFzQu
HtwkeSygTx/LLH0d4Z4xWhe2tyxzISbvUJn3vrdOr37zKoMyXrWBrUD1qEffRozgv5kSyjHg/RzT
qlpiyQ+qni9n0oPbL5n3WKl1ibnxAUNIwalUCXzsv8Syw0ekdIn2ewd4b+9XZsHQs+H2j6Sso5Qg
iz2uN2mTR89lIyMHGGXn6wHx5xZ58c7herSZiZRpS65FFmagOFhaAfqnxo7GoWNM88afSCJ11cvW
0J2dHw8CyiLLdAUMaFtaBgOB09djPiVAc8Bdw85+n/xPbRBDC30QmTtONfM8I9FdlJ+3F8ITxfQ+
RyetNNjJB2OFN8N17cU9v9OrgslBPfHvSDe7wNPqJa8aNS1noL2t7RNIwcDbPj4FEwnXmYGdbT1r
FJwcefUnVx08eGlq2QUOzgbO3c5+JRbKbBPe+HZ4piSYtXOZps894p0Cd726eibBEYsBr12nT/dS
7J04N9VsyD6iy+YbzaFu9hdlubFmhs+n1slsSBwe9Hp8usA5fZapel2uxTH8eLBvO3YPH+7SpHQd
nczBuYWEcDpsSDwf6tHoVBxnMfJ9+/QjziMDaKuL+6cqKlDJ36aVQiaDqZw97PB8QMosopx+8s5t
3WpeJ5o/ClglZGaI7LzTgnE0LrlL47xkMsXWgENJ+80IpCn/rJ/NZleIvuG6h/GtTpAUpjObMHxt
rVNGkSXcMwEBs6jvbCPhy7MrSRGtVJRvDsB69HA35WWpINCT/V3Hz4vjZYb3/GGoSjukBbNoWUhl
rpxCVmZvd/zc851aYehKKeWHAuKbulUVNyNWkgutmSAQXWEU3VqbZY/axqJ/qbkKOu0bclbP0ouk
4mZpYPwbLzbywg4iJECOTqdH+XTpRFBgjUXUxwYY+g6VHcFEUkdXWKsW52TLgCfCc1Cl2HLV5JjG
b4DFhEVu/cgRAn7iIl56rt2MSg0M1roS5wpOnWE4KF51eP2tAV0pXnbKISlrDGpxeuwpfTDpdhzZ
70+2NIiyoOr3IQgyXJb0dSUlGhSxbvQRJX470b2ozJ8e1gcOfpu8XjTpfbJClstoeJ/HWDOmy5nv
QnpTcPAYI47sxlcqm6O/DXJTWmYFYgIzyM/qCRrqcavQkLMnlT+dfbfyHihMScxLvO6Ucyw514wY
bldWH6MHGshkZ8hGPkXyyiE+FNsLTojL0hf51qK16zbA1xe/JKgQkhY+4m/O2zBjJgARKhF3oN/1
z2fiRKJ63JrFeihjZhWbWIj26ldgT8El1jNWJDkYIyRwkXjZie7nCViR9qPz2ebgVp3B0F948XFG
OQIsckWHMelA4OliG0F4Wq9Onqpoe4N5ZabD/Yoq6dRHefAcXahn8s7OgKJizbP64vyz0aR/rPea
NOrVZ2XAtremSSwgfaUBgh6I68kxxLXC547+CnIO/uAbKqJrJxUAHsZTkh08ofRKpg9edQ7HAH/f
peWUJv0+pXRHue0Qxj95S34/3Qfdl5CdQXFGPOouqRkuO7mj7OxABF3dL4d4FwMPKrXBslDQgNYH
01IXrPynDnLxxfQVGHEHt/hBgUoLMfFrqumaRLrTdo0W6xtzU2DiL3ug2aQFRMdcmGTnab2VfVcU
8uAkFr4ZT6ilgXyTcYdo1eYHh/BpE/QU7nTXkLMfhzkDVJ0hhFJEqYZSXUkZrtojdX3AZxAkqP4V
DsnCXi9WdltlOuPlP30p1wh5PCXGGYBt5fg6fT1uE+1Z4eBhzldZRzqlSljf5KBRajsH8K+HTZnJ
bGihkvBHNyKZikbFJ1NG+nuVZojouCecEyhe+oEO7HL9fLYTNLNnPZDAgZlUx9GhQlvnwlwiTnUq
RltmrhB++ucmi5BGWnpLT9I6fv/4hVUSFnoA5mn23frs3tXP70OTPzpxmSl+6LdjuR5cDn5k6+6T
Lrq3ch9iVAubDl4eUBoXZANOegCKkhXn2+3bTlsCxgGi9MI1K6KIE4r9Yg4vrO7c1tLwrzBPvpWC
o4QhzT5+IDNQYazxqD+0e0aLoxUMfJCDS2njT7lzCPipOdSoP4gV0s1ZiyMlLHwy4ymN9t3C7y06
ZhHI4g2Pd9Cs9EiLp7YqhQmF/eFrVs60dRTNou0dXqVhBnSDmCq123JbF5L3cn8jRXg7D4eDz6wH
hgfmIXDUxNN+EzaTgx+ll1RAsGvPS4ZPnBBycnsmT7jccy07WL0BJTLxwq+nKLzITAi/vXzlGNxo
ti2He6eRVcLklMDoeGDtBwR6f+bGvJ85nQkdYTL6huh6pm1CzrEL2YSOTdlw+w8z5C2s+5lfqg0a
yoB81M6iw8DRfGwJcZb21yyLRDMyyCLDUYnDjEbRxR0HBbipXcwm3GCUjmIdPEn8tdhbDlTqRcOt
ihC9p9mTSLRRWPnRPdoC41pEsH5oegii3hBsOyDJs/TTgt8G1RllEwehjY6BVjUUtBtjmeTIEPeW
yomoWtqXHF/RJyzD8Sf0eoBo6X+VwTXgS8HMXVZk43gKl/pelzN/N3hGO7lGbetcyzOqjUgVsd4S
hgtgGKDgD8BBBZ+E4waUWjaiN42Y78HO1a1az+BpVDruHDbo1IYPlTPrVVE8Own8wf63HrEipnvk
BqOk1NBSnVnd8eju8KncAACKtIjNesWalz8tzGyYC/CYmbIytzknN/OWYdeFpEAX7rRGMSlLWi4J
bu9F/wBcGiab8udHL9WuQd0EKlAQkhGc7udNzictOWZdr4BAVLCk+ghidwHJxWF5CFlgotuv202i
6J7Pe5kd1jZCHK/UUBIsntwurxTmGZCejxeZF7Up7upxKz/o28vdI3UJGAsjhS1N/k4isdvnvSPR
R5bP+R3FK4a/sPJBL2LBp6I4ul1GQ5zHWT/5J/LHGpATdvxTPi4YworB7wp2IECGLdPKu5sb/poV
0hqEtw7UbR2vezrI/xkstSZMblXhROGEDFeKEgWn2S9SzmK6QefVfvBK0cv7lbOjq68r0xEdSGgQ
hpYjg1nW/l780DOPDuL4xP9nLDSxMxGf199dpJwGdpfVa5HJCQ6s+TZHGUSFqEJ8KLR00UmpWPHF
pbc3HqTiII/6sWIs2FkKWhtcYZdSQkn7sgMZgUv3ZRWIhZTefr+Mwj8RVda+h0k2giT8oWqYVHOd
KginHxn6F+Ec/mj2LvuqT+8DlfmSS3TRiLNmXgoTbsNncZg2uDhosMCaeFrOOl9oINDkV185tncr
/9/+9YDgtSfZc8q2BHHQfQkNJc/HH487ctou67AZ1l5X+baev9jYtu/rQvNbfi5lLTxSDfJxYIvp
/wp/WKjUHKAyuVJaLU77jBclEVVJkjs/PGPiZAzufp+87jZHZzRNSscbbazJzVDXLSQexZhO2mxr
3sDyQ+v4lIwwNaMPIUk5yZet/3e0PYhhMcKCzj687ZWsNuP6YC3XpPjY3lRk1XW9jLSTZQTWOSwv
mZTCVDExARaxssJcVlWzPB6SUKWeOWWeoBkYPmUjn4FjGTMROgu2JdfWpaJ++thxWpDRW8vJTw/v
hAgmSlRWEIWvxn8iRpbiBToVbDMTdS1WvecJXEvNJfaBydxfqX2ZJOUAa99xr8TZVPOIPUpp38HT
uV4odXhmEIZ0rKAPFBFd2Mb1LMCg5PgE0VRtnQBZGmW21LTi41YlNNVAyj0QCElYRwT0cZa1uBhp
/yLvQNjkoOmycYaulFz2nJQAdbYKM0zOG+v4W+I+mSUfhi2shIEtUoMfMdURTjdoSYPNPsRztky5
/EE+GCjoWTHuyO6dXGBUmo2Bg0MKhvib1NxDy0JDwfXrRolUTaW7yPTVYHRhIuXczmo3L+uIErjU
1oOYSZS6OiTlvWwMmf6wk4t+qzOqErw97RCl0dL8wEnc2sOpi9z8xrcViIlgv818LV1s1ei3l4oI
Qs1Fz0fG5Jdzw8Tyjd2WCOzjDHN42yp7hfKwd+MDtlaL5o/D7CSgxCwWS6tc5mnD8goEHQ3VoaHE
UnfmzP/vIuFfS11FX9EcP8kxwP1A0gkyqu0609X4LRA9sTSROlF0EW564cIzgjUXpGLrI8wW43/y
2VEUxlSp6UoF9h8EStYUy4UDuP8trHY2x1MQH52ItbESN4xlkUFExjG/aEMmY+pHaoW4uFCVy1FU
PINElYY+WiJGeuxwsmschr73LqLKDF3jalLdgsaouwbEyGkzMET5cRJM+Vl87oSjuadhL++1h3jU
mzTIU9OW+Qobs8iHhMpAeGKpNZTMapaUGC75CdQ78gS/E3ra1+1zEYLFUqK/DWcOHnJV8Aet1cHs
y6V9E8nQmBKMzR7PVVI/e0RSxZwhtGfv9WctMWkJFM/aVbJxAgHHPzOVQdYGTi1IcCOfq5rBA9lR
Y6aVDvfn5yOZr3wInBMX0MieUnwysC1f/SdXRKLZ+eKL5kwgXT2B+R3CWMt4uNdBc/bT6V/XpZAc
TR8cZ6X671ClZhSPtsqIHLJlmRWzZ9kLHSZDvHyGm37aHRU8ne1j3zhJmdGjJ+gL8oc7ElZCZvG1
U/Z6XMaeiI+dODlqegycEWCyV2F/Zs6C3ADJW9dLLruMPSqTSpX1KZYIR1d8HXA2xCJuJ9uAWrTw
xgOF0WUHn2YIYlh/P2LpP2oWh+vgCiAd6JVUYs19CnAe8cuCnIApkEvlE+FiHFDmDi9jGXYQWUYi
8M9tUst3YmV4cFRy3jaEcXr5RCS3ILQZeTYyiEfZjceXbQ/11+3Et+kNlkLuQCS4qepYaXBSFvpw
3U95MFkXnExkAoq60Zpo7kPzoKaW7Sctuffiz2pV7UmFaivez19m/C91sabgYV1wTr5D6C8t4wDk
wEmsdF+JTgmsu/dcfgEpPx3VPCCvfWjEQSmvP3b0CcMbC+RPfe8aOowJ8QiWo7ejFDNNHzTD4d9F
J9eUUDkpIJqOjPz9J3Lb7Z/liZj/A84CKszAvTPNJz3Td3133DJJp87ChLmk16ACaIjkax34Bcfx
+LnawpkMHz4rz9qgpbKdiaTNEXAabwZ/sSOf4WIJYynUduzlYFOZWjRVhNu3L1v7Us8rQbqlaF9l
fmum+Y09yLxZrGpRv5QAZReUQDfVo6VQ3mQNpzDHvWVBgHFTdClTp2pIYZ+vQJ+gvPq+IH6C/WrB
nH9qNNVuGVnDX7ylA+cc0zDu/OZTE7eOGCyJHMMKp0j7BSlYQFI04z3Vpc9/+qznkbOkA324jNxo
wGfiIybzmx/iYezplkCWhcOrHQrtWXJtjNrk3Hsc+IrY4/2ES3KNCrD4x4LWLvZ5TC4ncNPcTY/j
eN6ZkvvaNGZrtAV7IEsCBUOLmP+va6s7zwclhS4q3KOMoa1yxGYIXEGgO2tjuxRDUp856LchMFCX
C4GF1C6MOv/v1f3mSZ4GYqN7q5j1FaXhP1vxgMYZRw68diXd/ve2DCLEwilZVS2XyVrrlhmOnIY9
iPHtXMMgnX0Ym4JKtO539H/S3bfABcm7YYRJKY5TDzAKvjMKZraDnSrU3eE51C6yTx/yU7V5aDbp
eNWRw4g/RlJlemcs02NxH1Wlb0caSLkbCoUCjhkLmQ+01G8b+/MAgD9MJZPsO4Snic8uPADtX5H4
6p2RLLonqbjboda3iBrk9pe1/Zqul4m2qOk7ytbNXZ34bNKXHbcNr2asFeQKLiFwtbBuOI/H/ucR
8xMxxHGa551oWQy9660mm+avzVGRP0T8ybaMy/LRnkOi+xkLaZZd/ZDGTLn+o4WB94uQOMfcjgpT
69r/3gckL1pQIQADdeR415JkUjyc/YNi6GFfJ974GZDDmGxPalnvHnxADLwVbPomO5km8PXEpPi8
RGCiLQj4EQJ1Jx42YbGZEsfKGKmLNCrAJ/fMHvBRm8E+WMqo3qH/LmXf16/E6emBq0hG2M4eE1qh
VLqQmsg6jGM2H5VwFDVDjcr5KrfdvBJAzP6qMdQaJSDGRTpUquRITvKXXebOFPdpV6V/9yKxbBGx
ViWo+jPk5eeTv2auuG8vylyrBXVJkb4DgGmKr9pZmGPtMo9DV/Az2LUtGbjCnwu71qaf/FPjOCK1
yH7gKeP3c6e/HAY5fS8j1QajTS9NbGnC/AsjHlXsbzkfUp36ljL6UHSqyWJP6tBEsEcaInOxr0AS
FnTAEKST0fPjPhbh1nuiekl2Q2vBtOnopKsbiysscitNs5YAOU1aN3ACRmTWSPxcmxGRtUOJsv9F
77fgaJUxAmONasVx/kQlVEuKpkHxFGLhyJKrhZ00XPWSaNTUSh0hAEks23zLuMC5Dgh0RHZnOO0l
zgAhgh2z7CQ2U0i13qIURbu3fNGPeH7w/i5lB2bN/uqOvXRXv6g3+UfpGlfl6YUyWGge4OwyBe+d
zmXrYqa+kOHNre+LwHam9q3pAcqT7onR7+olQfh7n9Z2skhxmFurQJ6FX/UhV9fbfm+V/+UDKi0B
A0vaNqwYeecdGHQAAghnL5tyOUmKj58lTCg2JnfUeQ2iVi4dslmVtVhimYDmcQmVY71/38FrUdma
aXkVUiskgKhTe0x4SGh6Q6Tj1t5EvO53CVZX7qq3+oILxWwpBanVqmtsGHcGzH8lEIutrJ3AaoxB
q3mKK3FVVjRQucYzpqpjA6SjjrqX+WLo5YuPNGH8UqwR1S/uEYsDaJLKJRAXbl5r/RhRtaT09wBd
skvTxmElg9Nv8LN56R37IuJ8C4ZWGtJ0UvbbRYNZSlhIM/GZWlzpK1ZkCuHyiiJg6iLv1ynewVF+
lJtRPkOuPB8wQPLZaT7LWCDbbRfp9BPboqXz3eP+7Bn2WshW1cAxvCUZltzrN4OdKAfBG9cgB4GA
A4yG9uqeRD9bEUZSWAXWSl55sJzJj6fq7tYFtE/ZyDRRYfZBuepvPj0kKn41vFObDQKbaTN1CjfB
LJYMek2E7hPQ69c2tiy9wY3wYSl4XyRvylcO7YUO4b1qMUBmJc0+CdrIQrhf/OQVb2wG/IqtoeVc
8ETtOhyyE558gr7grBgq4Y9K5O/MCTa5GoJpANT0FTO+BRnJ6LTzqdVhrRpXoYGlBIll3wEVLYwp
KjzAQ9jV+HuKk5dz8qsuK4fKs/EZBNVcTWtO0jl/4RVNl9M19E0PYSEo2yYGBhPBuwVDMBg/R/er
Efh99UegWFFHB3KO5vLyIJHyeHDzN6RUEEEKKhzVfRzty+t4qjbNLGfcym22s8ABfLyRGejrnRuN
5HfRh44dvBp/phbQCkeIogHwNAkaWNGSCPR1Q9ZwMtcBOfpmtRmFN/nR5muNUhwKO/6xRNRm1oIR
eaTtH3mGQG/JtPAm2BKicFG9/ilCRtV8MTqcYmBkSJLEJ/cGIONwZbM/zuHz2NqlvISW1CxCX8UJ
Q5H0n1SWWoNdcQPAhXYI++trmkiagkLXD1tcDIAyOLwQHW25lNLAIeWv5FsdDuGAoBGaPTr9eZCx
GkVKx2My9Q9Gwy5n5+JiVnasp+dkN00TlyOuYnJk4Zhn4hfvHmfit0wOGsWURJKUi8x8uDvkPxg/
+BFQntwFSX77hWEi4DHjoX6YOm8nL0G8V+0DzB0t4OkN6BNXClFei7SXjTPdmmj2kKgS2xJW/0xA
1f+qgN2cnV1N7xOudBrNBmRMIbnsB3gc3BmpamcdemxVQVORdDTlAncYTJDPmofpNTNCqhvNM7Wa
sTozb9pa2EYui34CKgxy/rWrtpweQbSkDJTkQSbEKZynrrYY16qLsowTNgk+m0atkl8byVYkVWKz
OAChKCT0402Moo/C/KrbF94SpyOc9UzL6+WH4dVDHBqRPjS/9bvVaSw45+Ev2QzVNgRLjWSVzeKo
07khp5AjAaNvf+eVP2UhKTwFalAleo8cuWGkjLkPvoJsBaq9/ZmZYXuBfYu6bkM3W0z/1bvWllST
b1/7rIAsxQ7ncnU9N7bteSUTdMYVYCE0bvtoYssV47t/3Xk0RiaS1XbdlnxAhANoTxNmEKWyRY/y
jwxFw1amTNAF8j15axMWbeOKam+gOHoZMCFeLI/Btw38jAqJpyu546dhQi6nUzHYdDndN21yWU8p
cY3xL8Ak3YcruQQ12o+JiUTsyDM+YN6hHqKvqzANJHVXqM+P0P484obnfhmJ9TqnXheCa7A3qO9P
vcq5OEbn+4XH37BMZWtTBw38s4506lymUURsWyKIpu1lxZMV35i9cEQoIh3KbmRyyeHub0EeTtH2
OpzXIZ/QJhuBMkTHfrByX9WMKYdSxtcwOXgTZPCkD7YUcNEPgQKANuCfYiJ6sHtVJis2VBBXYJjh
PMYPRZgK94wJRAGldqkcG3rTQXvu4lgs3hnuOg2FEb1VyAxWY5DB8/Liym2+XepfzxvVmGZHDTXr
mFQqLKp0Brqoou9g1/ET+NJbvc6UTEUxKcNPhTGck24Wf2SI4mRUph25guQwTYZ4DRJoazHFvBjF
pmCD2yf/lmIfXRTP1Tx/dkr9LDU/ry11gU1E+I6u4EnXbDp7PhwTC51GVNKqfRMvy/Xz+T4+AiDF
xXRIpQtIs0Rbf7WppWNDf+jasVwDuqxIBCdOZjdx58+1JHNrwdnGz5HtfY/FwO18TImaMKdu7+78
1iv0M82zd36QIpwoelSup2hZOsdDB+718bptOBBuP/tscyvSfBoEAtilH7iERNsfc0hUrEWy9BJ0
mbqGg4UDHzwmX9YsUoYEro5GIVD25mPyjQnQF7posWQrPtNwPlLuL7ouR5xBuC2wqltrEJeYNLtV
rHWik+muPRC2qOIi0jkrjQaI/ibUIXImjdEbYCYwepTdwWPrr/IkKCYFSbZMC2Cf9eFmcUUAJu73
2YowihBko48gFx8KsQLn45HCAnDj/4me3EpXGp4OU7d1vBNv6G2eh25kA3TZUKt5Gf4fJC5hKekP
gh0YA6cf/LsS8yaw8qVMn04TM++lPfn/pZadsm8t1Wz9nmcrLA2BHHyrNwpIZbMHIM3YpWKFaigs
fiZNX1GExSBjo/fVIRShjfKalRQ+Bw40KjE/ZKv3Wzj960DAVR7ySfn7Z1eB/Zzc1DNpeSuAPNUo
SO1IjqZ4dcgslo548aJjS3VPXM2G3Fx/A4/9xCkzra6ZqGyV0ajyqglCwy0sUnP6+G67rqxYvAqP
UiSHFZxaw2DTPpYWKeTbDgKA+noSJ36SAJYfOXABzOaPPD/gwIpuuOI0aZu9Q9mPc7Xz7B92KhNK
ZK3nWobXTSX2m9BjRzjh6g/7axhjnUmaCjG6wftvE8SjoAe5NqN5pYjwpGb55+w/JA4oBq7mbB9W
5iLlJX/UPjcAJLk9141rUsrreqWPaVJHlLfW7fogmHP2XV3NMJr7FxvghN0yu0vswwOwKM5W8ug7
p26H+mC6ZmMk7zQ2Hjct8kIgTZkpk282HCUUB7zduLb0ls8tNARKww+qOPasXQR7tXHRMwDpb/xV
c4HSP7tMjssPZPuYficqy82OIF3SooqSYQSNQTg6w5JwO2JrSN0GEBRIkqmJfFDW06FzIIdeumVZ
TfQ8B5tBoJzRtTggg7Z8mJZB28yjLIIUKgckk/yOBIq8oijEg4Zok/bOmF8WE9Vow5zWEks72l16
yC48v+Hw0gaZKe8S4RGWXoXwgC8SE3fpibolGn3Re4F/sinUyepv1bf1920nckAr5K/+PS7WT0oT
s/2GhTOdPCWLs/QYIOS1DlUhSBgfXYL8izyqZUXIU+IR4ecj1+QITmyLDzZMDUngHkuj3Im7NC6I
sI3rR7jFi67wT5UCaYls6WsBUzuug4VKdoEwADJJPxphRXmv2UqMugIoOZJeiOl504wKU4iUQra8
wQVn/yZUXpfJJc2IRxMPRYsucKy7WHYB2/7G8kU9PRmXN0nNKWXO3csp1aDL4d3ScHlVoSJM8Viv
DlpSFZJ4u2Gv/WKCtxDQFfhHhoPQmC6g4sTsLJCP0PQL//oJToeIyxHgjs32RiW4JAiHskDs4dTw
ZvHklDCAZ/5S1wnGcrOCKlveKRkaa6ZdABwOkN6ylLaSLmr4ANtKYz/vGGh2j2yQ0FdRvzaQ9GQh
bub0qoEacmrsvYNJaPFhsSIMwsHAyS3Om6l1oHOzw4m6AgJ6KN2eVhRnIC/3BkQ8JJE3GY2/0QbB
k2vCuPr6ItkpYo9Xj4aUnl1tXWPtlpbmJgJ/qbaw+K+jk2yrlOEMgPwzrVjK9kT4f6p+xMExlwlw
mVeewTcclC5kL1G1seZhjQgwFL90OlqPvpqtl5T8jBtPXUCF21x4WTFKuxoDCSm93H+qH1tJHSGP
LPUoP34+qqLbrugdWqqgH15e41eYBt8Jpd8ucVTgb0SdGGFZ5J9Vvm2PZiFsH/rGOYwpHPT3bkck
4dOTwvCV9gHqkobGFIzgP+LE1OSw7Biofia2vRmf8myy9u0M4dMNqn0nemJqXROElxfhw0VzIgm8
GoDJA7LAmTVz9q13e9tnc79SVZtfN1zWRcT+KiWW7S40Ufi66/5M0B4a1Yi6Mm2y5yooEAs8eK6C
DwvZ1ol4aU9KNDR+Fbf4fLuuSu2FE3H08pl40Xzl1vryZiWa1qJV4lKLShwz1m0jKz/jLcehIP3q
NV6tQRti4PHfXCC2xa/Vtn5IR3KV2aPui2lD4Rii57209g19J3sgCOhLXqI0Qlkrq/f2hbsItrhC
DjDsAP5aUwxnG+vjwfAs+7mJRqFeBiYvgcnJRbSI+MEdQ0ipmoUBvf5shsUNQtPz8ZisnbTOJIrW
y7KmT8C4xJne0ZSAZWUP3BGv0ah8XYznKh8otCs+W4l7v0ZEydvgge/ut9JQeY+s3VS9puwqdjBw
+fJgI3S5ZovKaXGKI7SR7/dvTuC8cBEyLDGxDQsqSROvfjhBCv0yVAfWiL5TtGNzIewcMgB7JFqD
PaQOYOCFfLgFK5OYCLN+Q7WLLfMT2CbsKME9HtVg+Xtjaea6ejXVqeIjDRrRpUczXdIo414ohPPq
hQ9v309Bw+WgFrwb784bNLpPkf7DAyKKJyuq9HYqlp+lhQN6LpWD4WSYcFPWCxmqyR+Sudx7EZIR
ZF9ib10xO3CEjQLFI7mU23B7fOXUz2+1GJ3U2pfz0KM0TP1HA1fFvq7jquvQnr+Qks2QcOluJidk
Ek74evxe0z3KWR25myblSH4ceBr6VYLMWhTMjMU0WHdPwjIFAj/Xix/j5bfZoRMiw/NeH5ePzLYq
xlW0ktbdnG1gzSnY9ds/r/0hdzp3eb0raTgdjB3qpQ0XXsaDANfZq+1eOxqpD5mPyOlWXx1GFVmU
CYw4ibKhMvU3HmBH382BJ7lPOyuh3I8ahmc2UbUuKXe7uy3dqmOYJxVhcvCUL8CMlc2tvfIf2U3w
vyNIAs6HhPsUFsWUvArfZPbc57zh3m3pPM/UQ283XQ4UVw/WAWluJwZPBbfJVVfvYfMi5au41Lj3
puZ+KFVe/nnEd8bTssgkS7RM7wXqPVX1XFZFlqyLde+x036xH0p2iOkm2efxtPX5Vy/UbTeHFXJe
DoToAWDoGvJFMbqZ6urSj9VID58egDOT25+UJsol6IhuSsbGYy6wHN4n7QYPWlL4EDN6V00dno0Q
WAnDakV0e+swaklz1eGXE6LWV7IBLKKE7l3DHmcyB3A7bUUXZpbRGL6IHMD4uZ095OtnBslJUYaw
9F1vFsg9xjV1tLqDlQtB80hY7uik+OUoUuDaM3ZKJDOkDXBOeCYk6MpQ26IqoAlgXA7zXylO0KgH
ZTtAcCvBJMtf3ivaT8Gb4V+oxNzwn3/fwzeXgOWSRfFT5IMCfjvE7tAjWogaBiie2xiLuM2/c3Yk
zv98nafShngGVvTNMIjJFqAarASFehDq8PxqzzJz3uC8sC44bVrINOl+NkjQvbo/pY03keOF+b0V
/UKJOzJRuGyz4XzSBYmewgd4y3MY0111UnAa7qMuFsf3FO5VY8R38OXUNB9jLDI1bm7gl6R2vzv4
siwCwJBN8VVCzVqbYfM69ZxMpH+bitwK6HapDGufA5KFvBzbWJg7N+adO9ZLhKHCxDATQtHpz0oP
k03943x2fOp7TXNwjEzG+c3Bp4dwP1aOgL8z0QCpxlBBI50yCLZIspSTX3hd8y4AGsGJFdyZhtHn
DKuzLq8CfAGiFbEzbS3hWn+FeU5W1OtcPOyGy433Og6DbvHBA6rmG7JA09z7DxA2eriDgeLjiHXs
XAH5PSqPf+7raQls3uNp60pbGZY2bxMPdNjvF0Vvdh6EHQAcXGaThXHSCOGJd6AwEdJR2XBtsVla
Enucf7+EmybXcXsZaBGTSWgQid/1qssx0qbFFQ4PaZqyEgiWOf891cNjoznCT8eC49Av+RJOoKVM
m7zWMpw3cxCRwdzmzC1fT6B8KzMNH37OJhwv1mm/v5Szs5CI+gEZtDe3PQR3Gqyk1r9wkSY7oUUQ
pkkKA6DSxXT8G58MFzyU2tlzP/9GR+BAilWo4UBh9irJREpwM/e+fbFkaVeii2/t+MoButKYYS+U
DuOhRxQPn9s7cDe+7r3/KUMn+3xLISl2QUOI4slmTKg+GF00NO6/gjsiBCOHpbsTG5uJdagRfcv3
QGLov97rFQKa3FudF4VM2zxYeLs+yFO11drTtq2Xyv/pQCPXwtu6UkxgoEqHmCWNMSTtRGOPQP8T
i120JDG3MtzzDjLlC33YtmuyzQYmYfpU46qoU0TxpqQMT0L4Zlc7Kp2LVuJGSj2TpAjqkay/7TB5
c9Zvh0e/58ReJ5UcUoKmVggnXs9nohqcjPBlt4wjPM0JkYa08PDQivU4AuOyuEHUQjvhglDM1XIJ
dOX95MPYznz/X2PVa5Idwb1opQpPms6qQB2jZ0M0AUfsifO3KAHBUu2ktqjewMcZXFL/d+uqFl4+
4z7uW3VWTE8B2LeQ+9pV9wxjdviowWGZwz6fJbrLXDr1QGm3jkC+qrVVn1hWUv97zFUp0f+Kcl5u
V2OsCrwV4oLiSrm3FCmO+0cQRt0VD13BhyT4z58wc80XhGgEWiJnisyKiNzBqHb7MA562KshXZ9g
WT7JxNkqkAw92X3V1bemxXA7ZAAzJpHtXvBtkWnFyvFkpqyO5y0XAXeO0w1E4ZxKIw9Qz/0hI8/6
5O9gZEztA6jOkvdbUMEEjNOFXQWBIuTxW4EUjoI3+1sEQtuZ8azYjEoiO1kCSj2EbBQFgIW6vbLS
/4rzq86HpRtnuptO5dpOMN4XCSdyc5CLipjprCSLC20vBHyNDcqiJUa1tkGbPlQVHhUSgeHRYF5F
j//4lNkECC3Je8H9sgg3S/X4lfqVxTsgOZm8hYG0bmEh+jdFZseXCKIsy9bbXrbPUPSd4lEO6x7o
djX6JqN8u2A1cFYrW1+EWZ544A1tf6jl3+RbtBhg8ZfmS8Z8xdwxLqrIOvCsT0siHHLtZ4gmOZ32
XWcrC3uT+yB5WOxPBIq8XUJecXIInZ0OcrRpoKsK2WnVVKRxWlcogbXVMDpB3v5cnsd8csx/rz1v
MCa4AVRKLmV26Rj9AvmmmLbme3na+JlpwfdtIYg/oSVdW7S9ugm076JgAM6oQea4JYjdNldWYQRQ
WRvog6sdSBd0jJ7IuDxkijpz+u99ZhAQmXEIjuHWoGJ4Of76jWvMtQ7qY2raYYrY0xLN/WsgmzMJ
Htkh26e5nuYykxKnfq3YcMAFTDvxq6Oz2RTQHMYjuK/eaLHTc+GwENY6WgldalfrKfnTfgP2QLUF
r2uzWHGfPdmeb4Kpxjewr13fMg5ZYcBeZvse3O+HFWVSNyITo0OiZ7zcEM51E2SFNhsnm22Zh25G
U25nNhtfGbUZzi82j2wZbjC2FkqE0UAdlfxZIRTCfG0Iwipj/fnrKu4OITHM92KNRgO265+Fvpyb
l5bQSS/dqoO5Y4MGKmZJZXjSQd83FrPf5mea3kpUXL0UGq3OvBHoxd6AS06mHT6EoTUZURr8aqhk
A/ts+f0ILW/o4+ZZrqfN1PznbPiaOT5+w07NH9sqoPXuJ2oaQjl9qo5ezUUCjyVcZIIWZ0fVJDuJ
/DGd9F4sNHJtCQ6qcfJSgWVMgkoO7ZariXChs/x8toUzaCrlzA8m3J8gGOx8mZvZfl/3EnVr6Fev
syUurA5HPq/t5Dr5ccYCo6IsTN1B+Us1uNWtBPxxZxlq6803gOqgj/Log0wdEEpzaz2YZxyQQhAB
iEcvlIkBCJye2tnPSDk837tFHe4bpsalyczImd9wELg44dEDQ5InscBYtLuyoPsyifli9t5INQKu
8sHLtvd1fN5Gz0C6CxVDL3rCPEzFJAi2o/Pp0oQc+Hzl3QDJzXu3AVcELklvmnAiwT4cqQaRYhpn
kTSWxnSKlezsCV4NhxGCZ68m8GNxc6eq1ZbuSDYgLi+V4DULiWKvPY8u4Q71d6u8467Jd8xWbNxm
Vre/imePZVSikm1iNhKHWo+z0aILD92ORadbq461/3/DOs5pKYO8fnz1NBLcDhqZVMdciwGu1enD
iuAthE4z5lu2pF3cbvf4hAohU1kF/xwUhJkSlGuBDAA8aB9B+GhrsAtuOwSLFIzMoALjpibZaQD0
aWJgvhcNl+4nWZsQEfcDn7YooHQ+jYzvokyayOXyhQ0zk1VWJ4MTV9zWcB2ZhkNhWYwZZI0Bkenc
NW2WlyAfruoS4kM9hK5uTDEjdS/0x+o0knffysFNdHVdWTtkexEeyvhQ+2AxyG5jK9MN69lPiVS9
HqCyIw3r+iXze93q/08SUt43ZVBrU2lF82QLgXahxZyJNrJ3pCOQqcofd5iVbzKcps/7kZi4BunG
zC39GhQjuvJxfULeEcQQwn0C6L/5XhPsvniwP3ezGfiWtiQmzRasTNmIT4Qb1pdkHczgdbp12jqF
53063jBK9yrWI3YdrcvtVQd7DQVX03/RnaF4EYtIcqD0RftAZEYZkv/jX3uF5N0RnjVHBGzi8nS+
3t7986+PMRckZTpR7GV0GOIfksEkOvcf5aesjS2HxawB7qcn79XQrjhnirtyNxAUIfiBJNIOBM0O
pUeU8HWAbrB51bTYvuc1eLf/y7Ezmlcgl7XWHdDx/cgLT7D4LgR6eISL89R4fD/33lKXpyM9zdS6
cLAQW+xkLxozlkMVBydghRKJgyLL6ltuJkJ/qF3ksPPokSBVpfq8hVXWxCEbPi2ONdf2x0JJOJJl
88D5HkdNHBs5jQissJAR18gKbYniLlA0bot0VxAnOVQNq5+eLQIZoIdqBNRTL5rwjVe32cS1N72p
aPVA4d6R6gMIc5eUg0ev3DE6xOrMZsj17G8ZnoBS03Oul1VPe6YvNYUgXZv92W/vCuJJdo+7A9nz
75Uy3y/zvFamdcFRxfid1Et+YuZOIZV2URhunm/VT/Rt4oSiT10Cw7Mlet/ib72V7dYTZkTw5lTZ
hprho6haRvwvtcWyFyChXLaVVTtDt+HSbbMNZVHt0bYZPY06QYW8/ZYnAW7yQ7FUjPQwqoafle/u
M99wU3lc9n4c31M+EpOZGeRzR40KH297eu/juWYYXa3vvZWJewR6ewYL8nmjvUoy4m1SIprCVsJN
qqnP5SPjQsbNl2AokN9Dc6IeCiN4Cwb1naMaVKMPVbYFWLz4ulOjDSEEa6heGKey+P6WmwT0UplW
mdFKsI2yGp4IPbk1RSW6lyGwqqThgtYsKQihR6WB+aiOxOL8BVCXO7Ns1Rarq/gXGOuyuRz1S2HQ
HoGkXLoRZCJJZyD3Sv0VDdOVa+ljuk1U025wf/byT/11dFDrxK4IlxMUoAx+LvsXsSPniqkOTzT+
uIbjLfvqIeBagWyIgTw0B2hGNC7qzHb6Mt3/Dr2W7TjYj4EAO/uDR7tZodZFAki38n6BJm5BRsaz
WpWrRnu7JGbm6XzfDHmNQLPyqzl/Lt0RsqcpSzxPlPwp/Qqm5c07ITOclbu2Z65DHmS1Jq3nQiOC
st3k7kCkUdCXuO6OPFxBOjfyL3q9mpJfS/5jGdvBbOkEJ6ayRG1nG/9WZefcNsPIbM69BX1+RgDK
SgwfFZS8X5ZALv2G4O6t4MIJbOm5SYL/V9ImXx4Gu6+uZi/n/aI8jV0vK2h1jfDXjDNZKhcbhGn7
vGFfi8cZMolghDCVF8V9fEd2oybXVZq/gK0IQ/205b4fZIK6VrF0eHB1lCynz6tM4PWHEVkgxSbZ
TgEbXJBdIXf+C5Xj6Bfc+CeRTOf8B/zPJnPc6FzQ96tNYKGM2in/7JPUPyxZ7FAjuYRL1SOHreLn
BSJXemohYVrFzHaNi+aItyFJCpuO4aJpfdcLoydi7r6FhaH1Dh7VZeqNE0b79nHaoHGgCAL58w91
WP/XXd8gzzPmEA3zq/5DkYJ4PvAlet5LdcB5/n+sCRorVoyPpniZi9JcMArv+lsAM1xMF8yZwu5E
nl5jXy27zo2K/sI9k0x4t+nPzRYNXgmdUoaWE/HEWNpPq7B9/ByJxX1XyrYbjFHbvM1cjTbHg3zs
KC0fN3JyC4+Wovri7F/qyzWBJgnU47nPOANzvvnJygflIONto0mAYzfACeNYKpPYKPpb8sy67VdF
f73mcL2KzsVM6tOED8M70DjQtE6lpD3/4VgZQ9f+8rW65ueqBLqR+PAoEwcqwKVIi/B2714MZD3L
0SYdN2BijndjBntgB67IWZOtBg3RmTHcXfzXurGQD6OEL8gwlSqzRBAh6uvDDkWHlvNpFOjSllAe
cr7ScCTVCcRyuuhZfEiMy0IpBdyK8ajTBxaLFaenDYBYgsztEmDq3CGw40cg8FmN1pHO7T6b1wSq
IkATpqBXell53U0f1k/pF+rIkplSIUKxJdaFq7FWIO7HPTyy0xDpZ/hDOfhWttfNmJXfRtOAHsC+
k0GQB7rloDFsgQxytEAaymdqxFKL86DDdnBzoeKa+4+RxsteMhEvbneuPEUfTBBEZXOf+DhO3AgW
Rx+rxNt9ZM1HnJmHkTcyruN6o/tL+ZwQ5zw6zHOE3ZTITwURyv7BhcepszM1ajkheOty1dcyCI+T
1YjWwyWYJsXQwqAxCDNYo7Vf5/LGgKEuRfvS8GwQiT6l7vvRwh3gqdAL7ns30AV1jZFSW8qpHctU
CBc6cfSrSTMa5w1vsFFs52MqascEY8E0crxlHCg64BFrYnM44RAKqeSeGG4fLquSre7JD4fw92sp
Vm18GJW235FAmqcgajnV/PLOEcM4s6IseEU7nD2QjwRma8HOztw5ohdVm/AAvWoG8ozsIFuZ/uoH
1AuY4ojFkVQ3rxZD3nDHVsMqSMo47eagLCU8Tqe+X2FudzMRTb/yXOxTPOl27eyRsJbKT5g1OiLT
e2FenPF7jYxsnbsmP4ehf2U3VEyzegssnM+8G8UvMLYlkSkyz+fwNrTGZccrNMqrURNFnKYtaGcr
/Nv/juwmOr97AogoI15N2QOOZZuvZ7ma5mWk1fiSZ7R23uaHVFu4x4Khf4vrYftQCbA2phTsGBLh
coIC9lB5DZWXhRuoVJIiQf18Pd59dxlFhanlTsxMGB3/uWKsizzwMs3XezKjCs5pfgei9gm928Kh
6o6C1kRUd0Rp7qKjhJrS5l8Y2z78pU5s3HP+YE4PR0PMs/WbNYdJFfYfdTHDKDzx8KYzH+pFv71c
Dc8I4lHyAQiLl+ts/jggYwUS2BSaLXnaHtpoTkvQk06b6xNaVQyiTKSkwvNU9qOmUG/2thB8bgEe
zn/NAsCj2mSParl/O9sKqDnJCuRAylaTVtSDhf2pQsW8ZbYnEqQM6zfqLBizyhu2W5pWGeVSAHpv
08h+20f4hy3JiPKpEnbJCZzHkvRk4v8nIs3GLeZ/FQCfHPhs/cIss42tbBmv7VnffRk1iseuNQJq
9OlR21ztADdif9Jn+0ORdtUqmMAK/qsH3fjU8Xy4/rq9fp+51/jj9vwLTgBk3w92DgdoFAdihV5n
uVfIy+xzkIt+PLh1AhDjf7+XNG2ifLbdJFHk+7K/iApj5wtDzNzEQdt2+OyAdc1/Hq37KJgqpyNY
EsfsevIXN85kJZfJ5PaWM5I71zIAdfZ1L3qbyp1/xVd2eWH9/jtywcku4locZ1BIUG5he1/Bhg0/
H4961yk9epBq7MS4OB2vCjmlNQg3v1hl6eXGAOw7iKHeTlWltCnHSzQdqR30ONitZe8V7eaxJ69T
Cypq5RAMjsEh8PFJt8inHcmLTpQ9WSzrzzUCmRzWKohVLyS4iGAvWXfJILRAaTXIEx1yBJsXPXwh
8iQNtxxYGQKb+0Xs91mjetVQ20F95Xs4HiVgSptV+14euGp/1AYsfd2VnvaxkS6t8TTho8H2n+tQ
LwMnypKafDLfIjrhunX8mnBURut+hyrUN77Vqa5DJcTV3do9QhHvOsaA8n3Mw/ndd+7mJhnwcD0W
E28KX71lfCn4sWu7jfL8jWu1n7nQQQb00fwee+Jx2Vh1iz0EA62/J93QV1Z1deBH3bj2cK/9FbTP
KcqraAwuge0ykNHkDrxkYt5t7X2nwDMeDAQpEkS3Qt5B/hcdWOvnRosQDcXaZJ+f1a9jQ9RnO4bY
4K+zSEKq9LHGY871TO7k9ZwPP03qzu6AiQxM81/Y+EW1ELkqpYZYvMUT0fsglry1TyW7LIc9XU7f
hOYasJwKGEaDbVHls15BogBU9LHElam0bu71Dn6DhJck8zQWDKlT3sP2j3HFxOnfJXei2tmmZt21
r2Cj9RPb/ZXSPpDCMdeOrM4dHPaDRrSpV0iyOBabEi0gUVBwTi26jjZMLJ47or6Rur0siXiQo+GJ
MpR2LarH3xdKV+SOSasdL5G2G3WDeeqi7+yu4LwAM6GfzpJGMK/NTaafRSqHLds5e6lITVi7ZXJX
u8pQL59h8yA8BcBVZmUd+16yPpgwAyJcA8yCCJmz4vpw7F/c4Xdi1VsaNfMy+KytUq/eza3ePN0v
/l0QMS0SYaSXfjIxylcYTNvOzgAs1yRYrgcrw66T4x8U4XcfBf08Gea6z2t7hy7lciyopVBMC6bX
Oqp4XxpTTacAUMXKHvsWDV71J4UQ/QoeitarGvw3aLDp1RWqitGo8KAyyMfsnUgYGrRop3pFI2iM
5LvrjrAO1fgINf7YXgb9bj/NuYTzGAgs22r996BhAMX1WrxTLwACcI8kOq1XnJUpD2eESfbznjuN
IRtFTs4/VvwYFKd4uvCcHHvzSEI/VLstwg9w5/JCRLf5KUQNULq0Q357sX3YcVV74YI7nJr/EOPb
11lCvvKt6gxorDddOT9v7dPEZX9Mnm/jokzSF82oZJpxlfTCvH8dQQsx0lt1TjPgFp4HRVMOFQc5
Gc5RULXo+a1D6AnvREoJ00ulor9Zw6ebr+2bxHH/jX2ATGjTJl2G7agdQXxEf0RV8U10/+/DgjJ9
jLwq8fVgqJ0aFQBZCJiEqaknkXfzm9YXL5i1ktLxvWO9MrDcMpODEUS7lj7xhg3Nr+zNO2dnarXU
q8N904YEbog/3ZHiPKmeuM4v29OeNuxq/Sij0Cs170FMpxOqH1SUILktstu+5iANPAEIPtNUN3V/
HSwXsxan8jmcPvvmjL/w1/l9vaaWGVR3pv5pmDuZjP2IyNY8grzPzoAQ/8bTOU0NNWFFMRO7fO5M
MNoER27Ixh/SIa35dw7fJKRsvuSKdoiq5duU14s0Kd/FUDJuqMuxAzNuFrSarh9JOtneOBlsAZBt
rZtTabwqd3ON9pfnLq70K7FcL2Qs2UM85gQ0FXIA3zCsaEaZnIUIPHoLE9EsgMJjXKI0AmI58MzV
CVcucYMdVJ7bjYSOQRcvIvM/KfNyNXh2e/Kgt0m7FRRWK+Vdi0q95NR8DTJ9RLiDzM2U/UqTjTVi
op0xggSwR/pMjRZEFaodtLuxBcgYzN7SePtgvLUmU77sUSyq2/ykbNNWeBbdx8crNgnYWLz9nSwj
3oFMSYq2nL/ixRhgKh+c3ERyxrytWRs9Gxqc6qpolGE3lVREPXKDFicvs231nnpaOnmVspSUwegc
1sgkJ5Xn0D8hK2YnkaZijNQM654rnwRgRYYHt8co0i1lxS4qW7T8RWIx6WKIM/zboCOX5U981zuU
Wf2xKo7KSq2GbehEsHEatTgO9v/OOCkuuMt+8+kDEsorP68mthgNAcwJim8pH+qVN95cZdnhx5iO
ETgq9OtusLRsnHe1lJ0Sw5kdbv8m8fJL33MeAAvQ0QF1+pqXOIGs5dJsNlEhxJ7lN4UudHB8I7fG
8e5e4NHX0Yf7TxPqise/BsVBQoVwUt7//cai0Jg4NZSqAItVelM+SjP+uuahfMYNucX+sAAVlq1/
7KKaF3RWg66l0ewesAeYjj59MT1WJhhe4tIs//V7H6LP8mXC1sjtmFPlkjeB0LvcscjBCRSKDO7r
OQ111zx/LpAwV3b03SOc2fiBn4qXIjH2c9b3aeGxpDtgb0yv6YCGrjAKW0LRIQpTlqexI/q8JnZv
nVQQsjlG7O6iiJhqwk4/cc9CfEOdxryVi1Y2bjXwzkvwfIFErtdUQPO2IOQnLgtLTrcZp9YEiyq5
oENVUgLBf3WRCs5WixEaGu5trOCxtc2MqSKrstQ8wOmiXhDbhPic/hBIq5HQ4BKyGaXH2yenbIHa
UCxK3tfLz7ORkaONbi2Mrha/hLelbbWx6RwBWLgI6vrlEcFqU1lpbrlZSOPmjbS02uAxUtQiWg/E
4EHFurukIep3Uo8OQlak3SwRAE5LWdowuKbVJ+3scXYb0cW7g+18kF9Zdtc3X96cAeofsEvL+1K2
m0usidiTnRUSt0FV7r9zfAF5hR39OZw2tr3p+9xAzIXls9V7YwfLSj4PdPuzrH491HAhw+hSsYyK
1XwwsDLN4kGMG0cwfNGZnyEYMxASblYiAM2obCYrK06mF9WKBG51n989e0EBov560WOzmkXSFrpG
jh5RT3ODnegLRbMGLa7p1xRv+417/gYNqNw6NBucTVS3mmXrlQoAccm9ksSvPHzKK1a+TYLm5D7G
Gx6nJLXNXs38Ll1TGLeqnRRuz0TORemTLWCaBVoShPaPFwhXzM9FxRzHhfLI8Owy93hxs1tTXZfY
W+BpCVQcWvNal1E1YpbSNKnm90osibjGZEnY9OTfvjqp8RrqV8Nrjrq4KewKmOobbsZkF5TSxvhR
EySLweyZN8WZibRO9C/2iT0KCzWs72dpLH7Ys79JfUSnwEe0ddinvIvl93fPKdoQ/cnCaUX8f2VH
hCsh/j7MZCh+Bdjc/3mZDBF7qQqz1G182k8Fmsrg0tTOO8OqqX22gzbs08BFLEXnhqAeFDvloORf
3UzOEZPQHft9HjPEg3NLllZ5dhHppMwx1IjCWLUvk3svrrVAeYqA2undIyz7SPF/xgn4byYMLN4M
FdkqA4L/D0w72lFVxTH4g506tU2QQjEDHI6ldgNhL23H2DCJNVdAXGvMX49S1/7vgRtkaUt0WSYG
0HwpNZh37CVOdI9UbVOMY7HJyFzMOsvxEZ58t1fpFkN8By9B5O3kkG2h2hxvS9jVbaSaCeWtMcN9
INdG5E32/JJtJQh3AJ3QagYqGtF9a7wZB2kBML2tK901vBBPI0yePgEPnHr/oWa3kbv0far8dKUz
axpx0V18aw5pGQWq6stxrEhqcaRtuj+RqdRmSNkt8Yl/MnSmvFvWU8uRtlMLu3FBSQ/0zB3SxLeu
A7Eq8lIddL48b562aBp06XQb1CP0/eALQnY6BbdGSxaXXNLb+gJW1jdWdckh7yLC5tsd+XR4lFLR
QVTTJ52gBx2HSq+JJhixcVD4GhCa64XstT0lkeOUxjCe3t/kjjxjv5fO5RxplfseYDhyCI9JEo8y
SUsX27NHiKwcf9+dVZl0qsMRScdUM1tx1s9cFJLbi6sxuldjiVm+DsB7lkdnnGiYKAr6wK0F6gHa
psIFGmCMVklfiT/ApKd8ACU5Va/mcEQ2N4ypzpOtpmotRGU5NIW3LT+VrP54rRXLtetn77ZP3Nv0
p/Hrr47yDhfXXfnYJOmFkjMqjaUJnPc5zpdyGTA9WZ5v1/zCXsVno2tVdaqS9zVSgrVahI4TqIa0
O75Qr9gktoxCSVCcjoY6FH9bUTT6iAhnrXpoQdxFkmvh91NVN5CdXLWo6bfcHsHhnG3PX2loVwMc
Vyup+MPek074tWyGaG461a7vBf76r0JqIYUg+1Vf8huRfscMA9H7HRXwOQJmGEnPH3mW8KpsLNJe
ovGNJUqM2N/Ng2Z4cpcq0SUpAXGHiGywvYkR7XS6EFT2vqXE0k9Kmr2GzFJpQ+9hftZzaFiSuG6x
314uYDrwgJxJXutPW2FAMvIidouz+NoYLbrd2pnssXNANDlfolOVPQW/aa8Yi7q8N5scnBgCX6RE
Gy2GtYAqGgNYHKIuaLreeQZCKJnBX7yP6lbRgq3yno4W4aWtB/HozoI4oUrM1TP4BiQDlHC9r0Fz
4dFIhmm771zf3N+Ri8YKC3A5b83p+XEMl+dlGDPxeTljA1ViDFCFVyORRV11H25x32P++CpK4qv1
uVZh+JxP2bEHrPVtujjUnxHc7SbK6bcSdfGkWZhziOuYhQDjgVAbeI3aNWRbnLfBZD4R2d9urju6
sw2ffe+QenVrGG4BcMSzFm0PTLZNSo1+JSOKjWo8KepJf0UNRCTQaz+EatzYMfE8PzToeXltyqQ+
Htx+o9sDzXReWEj0fDXb2FPJdDT0gh97Stz9OX6vFGbqoR60aOjnYzijJo5tzyHVMwyfymO5pK3E
eVoDEONGOCiTXK0/mxPNs5B3YwMXSQ568XSDT3qPjyDPMFGU9Td+WUfzsjjQrU/p44ZBBTNGdqER
2uOO6CcUx6v7PBKEbE680k8HZOcryu2kgmGwkRG5lbbmpSE/58AKCuD5PL7ndb+hjBGdClEeDCfs
5lfapljjAnVueF/JwhQ794FkpVEF3ziJ32tA/+VnHdod1b9O+Pqj4Dn1ccSYKiNuuMJ+m93E1iVc
f8ZLSZvC7s8YGwlyrWTSb6aa+TAjiVbTfwIRuJYiuVn/G0Z3Bkoe/0fekXA1gylcOM7oJxpE/CLS
uquFJlHxIYo6Wm/e1JBJWgMc1C4nncQK7bbJfwNGsHv4bgekMxeWysaU2CIFncNBZYGGEZO/Df7h
q+Q4WsckG35ynTViCohABNVvR63WQvUuQY86kYJN+yrDEh4Q4uw23ES5h3G0rm6Ez1taYvSmsy9A
lzLxyxefll64JTyCgicJvUUWrgS9FcZ47ZZTpCEQuhln5jKqJ+Zpd2bGI79RC9IIZW0K+crfw8gK
3SUTEeGDaKL4uNQl0XapFxcpzZ9ZCAfLIZFXl2hkkiOvKakfrSXk4Pn7LNdM0KouMpCkuFtSdVsf
9VgVULjZcuM5dJDgzRvcDu4uV6Z4C4IEg7pKDEgLorX6ab1UTnjOsuNAlQjwRDESr14qbbI1AOK3
ypb7OJEL2tuWkkz+R5ZwLR002Y+OkKC8bnK1E3COqHOdar33Q41j3eFVdZePcWt7rnnJTSUVFFzq
Du3Tq6ZsuO2HUQ1s0gXs/46B7QYTA1jyzNK7y0F/fC4vbIkDxNOZOVPQ5VisbTC1Bv5+CVuHEfG5
AXTd7xJSrWKaUZQ/5d3v5cWghv0D4L57x7ealeWXxw2trwW/GLoOK5r2Jk/e7hiVo45QzZNhfrXS
QYEnYVmx3fYGRwi4dDObDmkg1AuKmyF+a8JtX82j2NDz/ehuwxGEG/tW9WUBO0LPbSviPEzhsZuz
oG2kGX5HQqNSD7F1DXpufKIQLMwe1+/LPYA86WYNbnKvHV/t9T1D1mPT+BufSWHb9grlp4rAf+g3
bqKPHXc+RmtYazCPltiuWfavNd0m+6kYxa7aGIP20cO6Pbz8Z3sjoCz4wPdJqUHiN1pQETSzeq7p
/bdVGAsXYWVpaFRNq9dE4049JKFtiXbPqeFdW9d1gVCrNHyy4SPNn8HzUuW92+GREtid2gliNIIN
7q9Lvp0gLeVkBtOAlJQJblYInMkXLQKptAEoL1FII0wLGeYQB6fPRjaMom4RJ5BRrijKudfUo11g
+5PFoSKheapx55UIEFxJUCH63HLJMMYFnWRvOqqkOpNPxf4boQaQXrUZK/DaJTJ2JK0ZAJtyDobK
xZRN7ml/nS5SIpYn/2R+iJ9vgSP1VZOB353aZ48dQLQI5nAUyrKrYMdhO0OzgI/Ir+8dNgYY8Vuk
5MUuNRPiMYTt8MD0ZfOnVkmMxG7DhoagPzfB1X3YS1gT0kaiz7sRJdhwrOzEqNnVV8BqyfypbaMU
xaIv+2nVv+/FDM4J38LtMLCtfnV6ojb0sz0LdWK1k03NOyDMRtnJ7euORmvbVdC4wGp7SFP6PWCW
4uyt5ZwcFXg3VtbazBM/9LE969Yiqlq683vqM8glxP+gt3XgQLMvzUGJ26TFYr7xUBid6vu6G5sW
TlqtrBPX5PQJFCruOBwM0v1ZWiGfAwFw6uQ/gqKkIzNu6D8GFAaM3pQocvO8Un2njZWNxPusHULp
ddobeNtK9b8feyB5zRFHJaNHFp9khUWjibf64jOrd3e3E6koR3jWzsIhvvxRw48o9hcoQpzak91i
TxHXrtihnIfekfaSIQT+j9Y1IqhBb+teq1sWe57u5bXVGu4iyOLsFeRdAMXboArV9mU1WgqYvKUa
sMypYuZ1G38u9+6cHRe95n5PCwx9h73t4HhwU+uAQ/7lpACeqg0RY/3HjT8IbQ4yWZucJ2mNxdor
fJyXccv59LIAaDPRkTLLEF5UsLNsuy1WypBdBvemQPCfOMbnRC8sqpHQSWE7lPFg14CXlucI9nRJ
oPyOJ0YvRP8VfssSyZT2968w3Iz8bIE7Jl0OUlVh5I2jPqrDSNf8kWEgDaK5o6dwsby0H1L24M+J
wRP7xpH5v5DD9MJ1eWAuXJC9ejEFqbNP/xA+bK20JxQKHKIxzEKzVvpdn3tXqVd1tMY/AnDB8Z/e
f18qfKhPLNwD9yJPMq0vfscN27GlQwbvGlByG3UVD99uzmu4YMztpDjVKToXrmfcrnAhSKfwCP8f
wO8AuKswiMMqs+RX/2qpAJFjjtqg1LO5vR5bAxiJONukDrpKm8a2iXkbp3IR+MTqoetLqhCCX6Fu
pxoO/0YBYRNECCLmy7k7kCFy0qlGPMiSiqSNby+/FREOkoyOLE4JIWXZmtTWFi3Zv1UccK9vE003
NrcxjnF1uYRhzvRZHtoodDjp9+f7eKcZeljS9DLCROf4SHXceZ2Rdl6sDJOyZOBew7NF0OBWb/oa
eUsVRfzSMC0Tl/3lZtVLik3i3TWCQ3aFtQKQ8k4dRYSKUM3vOVSDLN/EQD9m94W2PbUeEPYsSJ3Z
OD73hiP4F2I98mQDGHr5hkH1ostbsi3lQ0bImFc4Qd8kQ9hqZndBX8H6yevT+L4KzlqxvGAG5mRW
SP55UK/OeL7z1c98J0elCh35h2BZALfdLwUTxlBtQTz3zc/WLoUVX5gcpbhs/ez1C3uemTyaRZNC
N6rhPDrcw43LPoUL7NueHM3ZEjxFASfUMueLPkremvMVpruEpMSROWxyOetaqhBpCwinzyOtctOU
24NxXkWjX6yWlb6Jf8JujSsadfk8f6NQpOhqnybwfFMkdf9yUBYkwRkX2/SCBLSozVyLWK8nYLNd
zCQxdd0hduDz0eHgInf0mtmmIhV9aCCoBUAgJeaY3K/zeYEPXijL1q6FR6ByiHRTBTZkf0a18vZ5
USqwww5668KSqaZguyOXaimq69r2n89RTGDOw65IJGI1jpyxJIPr3z111g7vIc6celGpRHph2F2I
NvxuDSokloRJLlk+01R24ZXLnAa9yJof7XbAmAsJJ6dYBVIkNhGAuYEZA4DuJ1/IjQrVOj+7Dfm1
0Zpc18FDvjmHYKnpX6GJnwnYstmy28D6e1BMY5/KoPd36cMGtB3ZGEkDVcceySEaR+j3I/Wo6tac
MdVdHhoflK49MCrM9lq4emhHddQ7Hp633Uw0v2KmeXzq020hw7U94gTFZoUPkIO07r660lrTHKNy
c7BqWbh3mGQfB4ASYPLUYTETl9mJxRXtgLKR3yKei+ESkMgGsk5Zvx9Xrdt1HF0CSNXTS4tp3xCP
XFKY/FP4RqVUkaP+E1arVVUAbGx5LY2edmKO5uSBSgsakidWr0OdpE+H9j3IaXJxxIWwGSNH2D0H
A9UCey+h4H0ewcR3FFzJlGy+Zw60MD+amhOqNPinCBVm10b0NZnmo9GWK567xkvMskFoYcj9v6XE
pw1H0c3nx1Xj01QgWsTHg31g6KdOm4pgbsAfFg827zbhQ86GQweonVtD66PIqyncfJIRaENT6wru
yQURwgQSHc6LzmlKqEvDwAPt86ypcywtPHUO1+jHYj2N1muNw2oi1kt2/mKsvd1KQ9HpIKGfEnSR
+Wczai2N7UhHRkE4eD8JvBJHiy2rpG9QCzPh0cKmRiM7vU9cAxrAeJsTZLsslVGQzIQgLJawrn2x
UYdl9+bZxmLjCFQK69GMCYWYKLgNANVsHG6gHmLPLSJRqRv2L9ULTAj8R1/devFHophJczSSxqsP
YnmRLbgpeqOHOM33mfjuphpN4fWkJI5BXvo9TOKucGgSc+AWzda6VXZr7Qti60T7nVHeRESKyCdH
trWZVa7lG/5H0NdoY0gl3ieEXyxWl/FN+cc+lo/F5w/wv6fuCaODrk8SFzZ2vDJAZuBYEm1TLDDl
YRPyLp3fwdpOmtz7NCH0ZMxK7amwcvDIpkl4nmxPNvRz+B49bVVCfe6Yvq8ZdA6kOOcpA6nXCirV
T4k00ETekno7x2JHPy99utmi0Xg1OHsQSAVd1Lh+GWy+udGiAbt1YxAI4H0otn/I8CoMXtaqPvRt
bphwUQMLMpihpW1Rd1FqxB0sBpKvISjgF93K64yz193JC99yrxaCtOs+a5RmBMOPDjHzKToigS+b
l+T3kI30WxcJsNsW/sSeTIgnjXc3BZ6qxqvQWUjt+aYoKBAYfBvtBlNTLj3s3ZQr6YPraKih/Rsu
NJkCU0Pd0HwGsWCp5AExuMtVjM7ljGVFF483FnmvMBJh5sHbk8IrQjLsvws4dxZowM4/Q/m6sEYH
qYfpanO8BLcnk+9Hcc5barJtnAuVwC+bVrXGn8vgXNXCg7mZPz3tu1gzSulreKvRUMUl//foKZW1
fQrJE5YWGB0zUoDBGxxA04TrrkBo4q9Rg4D6CdMKMYdOgXFXeni/EgVaBu8c4s18kIaDHKFt7/OX
OC4CjHk1HBjWUVwDWBEgPAMHrpBgyewBrkh5FbzyPhTTuVNmGAqWqXw6M+BJWS1TKbIUArIByeTA
39hL8mVXTO8uCuB+LdaqaNCIrYKoQJ/ijAD3EvGkaOHOY5v6227CMToyu4+BqdzBrlGc7UnauCIO
/F2+s86msHrKc6t8dlvaPtt5y8fPkbQ6jzcXXI7/ptDfS4HsLKCOkzV11Mkr4keswDPd2zzaZFfp
AyqPdG/ZUfOA7yK2teq8c5lDvZrjeE1f8PjzRTVLWC5WTr0ZLY2pHxsD0xq0Sbpomdxq/HfbkMHA
dnJd5EfXStQh4waD8o2Zn1qoSdVaK1F0AUvFfDDZvUCKznWymfoYuWsvDea8YCpUecIgencHjDBb
NRCz2QhkGEMskITH5n6JYiVXRUxNjbTnpomJqcmm2bfRg4VP6/Fepr11+OOp0+AbnYBe8H56eGea
KRouEJrNg/2MKNLAztDSkEN7bPDSpotWkBWlqeLt/HP3yStcJu2C3Wo33RDBXMvlMOokh1JiMj4c
UZz7p7tpH5KPRT50Hc1xcOglhr9A1LxS4PXQiG1xKb8k3CzOrwprS7b0+I2uHt31MMTe/CxwRANo
vvpd9Eu7wcwjf1I47VYK8WN4162fnvy9uIZeYjpUW5lMh6glj9Z7KfvymF6zHgNB+YR6d+8rxPjX
8TFYKifhNmvNCVPDv2KTmCo3qsoL5wcGd9mm+0HKQCgHDEwtc8/TTkpIYTREWuWztmP3B7EZwHWk
gXz+zCviDTe0IHYFz9xaT8P+DaCHRxIkOS1BXJjy6ymlQOqQ1TnISfzFlbK/E8FVs0xnN2J7Q9b5
HRLStYqG5w9M9Fd+Z5Tg2sIoreIze8FxRbsrQ7LTe8MXjkFXsDlgwD4KFYrQKyNcpoQ9LCbB1i1x
vR+9a7KSVU6Fjeyff5biJFiue9FSrM9tWn+Pm4JV119rIqYG64ajf2+08gIOokG3lVlOLWlyiLGC
GOKXPRcEVVv0GJQ0FCgUbLVdzCSwkNaJ8THHmGfkcjbdhHeSrAKC+HmTqV7PrRYWxrOOgYYy/+la
Se7x4qsz3BwE+/qpnHXtqDPXIMbIsy1i3QU+y5l5jxw2znJCPCVH7gGmO6bwfXMNHpCdxCxqI3eB
28qogNUOQjrcVgAZuPqvLZBJdTD33iNxzmp7beeqDSwEifWE5iy5bstyGdxzSBUNpGiQQKa3IjFk
Hpuop6SmBNy82IQAXehpFwsSaYFE/XQSDjOrKhxNYrjQ6I7pFSMSg3DHqBDmxMCOBVMu52fepEHK
X5lcyiKZYusOzFuwLETDJj25Y05Tf0CegxPLvKZa41qJnllFVMVfknejz+ruPOIxpeOa1j9c3rfO
OVYJD4oHAxtYRr7MwgD8Ysj3rX1uQfBClIEqbfM3HAr5QhSaHyAz1UxE9/wjh2+Bz0GMj5V8HhT5
iXTI5vU3uFVaZCPqZ/BPhjyLWmdUSUNbWQip0yP/TRPhZS7EX2GjtDjRjuIWYlLKk9qXv2wzkX2A
r8+jewS0rkAx8t0GCgIpgxvOusWkAyGsAzaasyZ1M9xXI8rR7l7cXV75B2i/hb70S7ioTcDSrP6l
u7ymA9svcwQ8YhJEGRJB5J2kLU9+Vl7ibPfDWSAhwgoECw7Rokc/pGnUQdkawzsEzCwHuZkmaSV1
I9XbWZaMJDQTU0rQOAeI7WqNFgfeqk34VfRpCG2C0uL3PDQ9ktuNF27+o2w5HHuCWCDEIu0Kul61
dnokWd7J/ccwZ+ugUiBCqCSfuyzQO139nGgZcb++UTZ7g5EI44Js0uWksFzDBivjR6lRQ+3fqmj1
rkWjrrLUP0wVJ7Nq7sNFmZ7tjOnYajNwp0RM45vfetxlftxc5z7XL3BlfZOtSE1OAVmn+UJ5imjq
K7ATTKPwHDTH8v2FV3tFjBoY4m7iD347AQ8eGDn3V+wJv7mgbvM9Cj+DDdpXL2zVB5FQwwZJ8+8b
Wa+0YbrI+Pohg08cagw6JP4ACPeg/3Sh2AIA0pcprsJeVa2HzRj3TLhyPAwHBuDzBau36PPrdXEu
fDy0NcyD6EURwEUmcCEFAsD1cBBrk3LlZ+UMCrBWwY5hA4805Xwm9o0tZbRL3cAc+bTpRk4PNCuB
4w5tmeYhCNfMDoWoiVBCpmME/eFQRqxnqMeA5RBGRGHZKQOxObljy5LMYkuo19OAelVouIQvttcp
OAKfomI/tP39e+0vDOt8uMne6nPEsxY8AMhmzCm4sBLbpXZN5ZyvNpi63rOoBmKM7ERbkd6l2fxY
HDZ5vlW4mvg3oLz2u4vJOs+zO8Yoy6pFRVHhqJxalXQ3Rg7ZizQUQesCr8g01sSgywU/kdtqbJAU
PIBjav59B5t/tTS6W1EgP6XgFt1agpbwHPyqGBmWsJcnEeAoV4Y6TqWEjPq8Sgz7alO4UEZLw2On
+CErdLFKYbWZS87sY+uTDeXXvrOriPgSYAHQDZzD75UyK/VJvM69Qip63hhMUWAXRf3gkDPZHyce
i21zgI+O4i2y5Rd0C+L8E9+nNPLwekwEbH3HW5s9EDHx/oZ/Np7a7/4qM2zaN76IDqhZSNNbUlYG
WxV8Foqwp0ddhpIVBBApjVFkkucUXRrOvxbuUhhkuHl3mDvI3LjAx4GboXdVRdMDhNY+nxMz72Sr
4OFoJypPWNdlLH05/AuITKuEZrMNljehoK/Fb1NSdaZfAdfEdWOJFE1iJwvrsoBtn5GyQc/PqfFc
qcZhyi32Ne0IeN3Ev/oWmx6DSAOqDcA22jXjkrDH6Qx6T/rjAK6m29tWrzF5Cwx8ysYnlTyPiJRN
LrrRt2k5E0iM7U+6qu+N9SzzGO6q1JgFIxF5GmLcjjfbHY5DgYhkdnenZeOIpJmLXAehmIYwzUpa
ZQLK4qaativXm432OZcJcXiGIydCw0zkHPuNEpZPg93g65ww1klGw5Jlb/u8FiIaPqyIJa8yVGBQ
pgnw+Vc38wyA+7cDNiQLpS/Po9BPJY4JWWOhxXWmfNPXx6lPI6XqHPpaGtYTy7zALPh6VsQIaPWM
M2L2/ghOBwNAB0qZJrJVi+rsT9HQdqQLaPFCf8tdFvVZ2jIhtgKOAu3Ee2ZFKLEBuGjQ7MO+WJ9x
z15SluYclHMUJQ7yLyE9VPkhOVguXvIG4teJyYpzN6U4s43JCyJ9BUuxRnIGNGDOUqzu6K49RrkR
FnNTVfdKUjHlvFDLCqdkwX7NhRD8JGhQv72qeSZ6IPiylQOiWASE5wvSeHYQaRni2UnQe03pg+EL
aLsEl5A1UaL0gCxvkWrrCW4si52/DXfFq3L9Ta0PvgF4+DoSQmQ0zuXKTVGZP9N23U3IEqgbg+dD
xpa9ozVmtm96FE3+bUF8Oy56gQol28B8Aq6/egcw3KPDbw0MCfmuQ2w6ZpHfxQGvk1238zgfgKxb
p1SCBB/XGkK0hXthVxcjAjXWM8JcNFMY47YghPEkl9AeZGsVu1XZUfR916ZNV0njvtmhc/R99CbB
YdevWH/fOJ6C3i7nrJq7CgDsg/juQAP9bAwQ3RR1Kdco6Pqs3pHSSo0KSUkfrPq3bE6zvPIoorBZ
U9eNemfT4hcSsjjGsrLfHw9Tkz1Uk5d0cORdt9cVrUUAcZeE0+OdDd6vjol1UbgwBP/o/6yn1HbN
FlJztvjHnXKKQVeda9vEznDPIv3Q/b4EGj55i6XLZ4xvJ0bw6DW5jDLpnYtxdOM6B6IMnIMxpEzH
Nj1QwkkWdlx1Vvs6vXq19c3iQc2oNp2fr1xCgTNjG1My02Per6WfhHuSm7YBRChBdBefwmYQyaI4
JJS6r6vFp3dSTuTyscEn6ZzuPWqOlBlQfPTlq7n5WtxLlM/Wtx2h/daKAOSkfCY3ZCjnXOPsCZdn
je5B8HdH6RqjSb4AQ+kJ2plo7q/ZIj/S0KafxJMkD/CfHITKuJYWnzKupPMau0HtRSLBkuOYHsN+
BYQT7J8FFMFLHAHFY1kD0UDRlATgiF9EA05n3z5fwF5NjkGeJ3dLN704oEaC0So7FLa2kbY9wilY
8IpWv2dEfNQXMApZJ9M9FXQ1L0HJbVIzW9+X+2hVFiDC/NEb9HD97ZCKRWzf2uXN5tfiLfmOesNR
JPsBFqfKiXQxClRUc5kGYImsFD14gfu2OuwIKxpYxmrWlYyeS4ICLbbkeTekaSISLHfiVvzushK3
LotJLL2TvsPZVonPzA7dtBfCIEBj+uNkcW6mWct68PErWt2jt0VeRpyiJ3i/78FfncFUI5PiuF+r
4kmO4R146iq4NgapvhP2v6d3Kdkg8YiT7/xqRh0vMoppFuQv7C4SuqnJGzbwWN31Fh9OgKv+mK5U
EFl1mocsgog03JN4hqDA44wyUVlo5ImXg96jMYmk+56v4sNDuP8fhjXh5OV84SyGtyLykIJa0Veu
ipHmN2k35qk3op9V8dsshf7DGxf2iRypkP4j8a9atwa3mMh0uzdRw5XutVbfZcqgtalw1n+cdXYt
ks9QkNBT+8ElZImyH/8QvwL56tjT+e6Gc2Nsu69w/4IAUKL7M86FLlykjJLFDbd6UNSOtN4VksTk
/+RohFVuJq+Yj95DZjLDhM5lAtinAMtd6ylhYB07EZnOU/tYkVQM0EhPs3PDN/9B12WS7Sq4o4xj
lyqYH1A1aNh6C7hC4sTunhtINFWMZoOyQ6J9WUaliSReLnYR25DvFtUJAtTprVkStvb7p2sLkcxE
UEoFTloxt7v5mCdprv3RoJn8uih5+y7gYuwat2ErITRoIUCyjhYfTpPzUgRxh88r728ool1u70Uk
czTpJlOnpnywfO4lJYAMqQhzygvdLoiJeykzvdCFdd6CxISn+LpSkVDtxeZjgfkRqpekctn64xkN
+wQUe1tK22CbZYSvKQ9waDmjO3pF9cPzRlMty8i0aiwhGnXGwtCx36zME/bTzvTHxTabVCoV5DX1
/02OLbBsUP3syDanABKWfzrQneTc06m7Pjw0vx9wuh5i3Y3OE3O8mPnvi3qt15SeevaNwUTzTI9X
y+ywZzx/g3Bbq5O8aYDlJmao4TriLinVGXQXfrgqB+SwGdE3QZtLuEpVdt0LUZ3lW+/pUTttxaUE
7OTrDOtJ4vC8hSIkZzeb
`pragma protect end_protected
